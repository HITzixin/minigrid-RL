�]q (cjoblib.numpy_pickle
NumpyArrayWrapper
q)�q}q(X   subclassqcnumpy
ndarray
qX   shapeq(KKKKtqX   orderqX   Cq	X   dtypeq
cnumpy
dtype
qX   f4qK K�qRq(KX   <qNNNJ����J����K tqbX
   allow_mmapq�ub��]>��'>̍�=�m�>�-?�]8�@�Q۾/����5%?Qb>8�*��g��oN=-e ��/������sA>毰���>�:6� yF?	����/=��߽��>ɍ�~�B�zb�>tl8�(a����=}����!��H+��
x�;�p�>�4��o�>�Xc��	?�������ǾX�Q?ș���ὨK{���=ŏ�{q����=y�����:& �>���>�d*��G¾/vD>B_�w�8��2��ӈ����>�l��P�����>[y[>�? Y��������>�,x�
T��ɼ����>�A�=�/>�`P=|�?�%�>=.M�O"?�4�>D~���E�>>�2�x�)?�u?$Sy�im�=�"���^e=��?�o��_�������=H�3>���>	�
���d=UX	>�پF	�>[E���>�ˣ��n����{>���>ޝ8?�W��؛i?z]�=n����4�,�ֽ������=R���������=/����J>��=ё�>}�m�ɟ�>#$=yr>*%>��+�nRf>`9��@>Jp�b��>���>�%�r�?�K���?ͱ>���-Z��r ��3�����>���=�w/��B�>&��=b�Z�Q�k?J>FW&:��������*��ش���f>�<�}�4������+��M$>-?sn�>k}(?6�F�[W�֨�=%��������=��~���	�=M�S�n۽�u�<�G¾���=��<>D�?�zM�BSf���1��J!�V��>�Ԫ�h)�q}q(hhh(KKKKtqhh	h
hh�ub���7�;·�s����8�����D8�x�7I����7@��3$d�8�	�SC�54��7{�E8f�8h)�q}q(hhh(KKKK tqhh	h
hh�ub:�»tĕ>Æ>�݌�Ml�ŉs���>=��=��:�1��>�t�>�=��>�>y���&�%���Vѽ�[���n�=�-�gg�=G
=U�������)]�cP:�@�H��8=�"��Ӣ���wT>�n^�?��=���>mx=>w�y>"�_��b�1x[>~hO>�F�haF�U ^�f�r��H�>��Ͼvm=�W>�>��]���>,����=ͣ���m�p$�+*>=jѼS���
o���=&���oЛ��Ѕ: }���=�I��eƽ|2+>����%�V=F�>�H;��Mq>G�<�>��^>h�^>�7>- ��c�$��w�=c9}>$��>�ý}�u
&=�bm�}�0>8��>l���� �=�<!�t��Xｃ� >J|ݽU�(�~:���Ǔ��Kc��O���L�=>+�=��/�0��=9<�=�.�ِv�{"���(l�؉�v<��>�� ��`����J>�>��Q��=2'�=����3#���0�=,'�>mJF��B�}¯=��E���'>o�<�E�=��>x��>IY]�	���t@�>(:=�������w�Z���
���<���>�ɾ�l�=8�>q�����W;�>I.��1�>��>��=9�>���=?�=ha>�z6�*��܅>$9E�S���?*�'�꽒{��w!��4��FG�0��=*[r>N,��B^@�� �?�>eٷ=D��<"��<>[����v�9*X�����0>}�v>�ӂ>�I��=��=�4�>�=d>��C�b?	>I���,Խ��H=BC�����W�;7�r=�1;���b�G�h��?��=a�ؽ�>���a�=[�#>�}�>ڨ��I0��E�=�+,�3�>�騽a<�m�:� o��2�� ��Ѹ��ק}�&�/�b!�=܀!=����m�<>*f����>m��=�ڄ=�٧� �>�`=_w��`?���>�����>&�����=*M4��Np�v�=�R��`<=���w�P>=KQ>��s�p��=�~�=%�q��Xj>��<���<�yD>���=�vѽA|�ߙ>q/��* ��ʑ8>��l�Ϩm�8�->��#�P>3�W=�;o>�c?>ǂY=,Q�E>h=�M�(�_�9W��1�>T����U��V���y4>�A�:�Z5>��=���=e��>X('>�*;>�E=h>����^��=�}�:�Z8�[�=�&�5��T�I=`�����2b=�!��~�9>T},�ې��2���|=����j��ؔ��w>{��<��$=)x��2����A�� 	��p�<�u9<�8��׺�>U����=4��:$;�C �>�����>�E�Oҗ<-�I����i齃
��Y�i��8_�(�=�9�ne׽Ͷ8>D��"0�;
��=�!=���=���<�t�Wc��5�>i����=�>�(M����=��;�!z=.����d
>��,>��`>zO��ͽ�{a<���= (>
�3>��s��JC��(M��[2>忍���(!#��G�;%��=!��<r�>B���M��ř6>
6S��l�=fy<l_N>,��Zꜽ~ݮ=�>�Y%>'>,�h��U�=�d>��L>F88�C{�=P7O=�����$>�;$��8�ت���o�ܲ�<�n�T�z�u��=WL�<���Zg
��Aj�3.;�ׄ����t̖� ⢽Oc�<+�9��>oXj����</	s=����P5l>l;��>;���%;ӽN�G�提��>�/Ͼ�,�>qڽȼ�=Ew�J�>�����=���<��>�4�>�Qӽ�'l���9���o�ѯ<>9^��=ݕ� �=v���bf�������=�7�	<��nS��&�>��s��t�=o�@=��X>�ё>�i}=շ=r#Y>��'>hs߽���\-2>�C��B��<��g���=�$����=<׽��=���=>��=��>��<-[�����,����8�>}�>k��<��>��F�R=B�O���i�邶>�+�=n"�х�<ܗ��*����=`�0�<
¾dJ��!v��d�=���=$G>�K��!���	����.�պcĦ=[�ݽ�6�^6y������{N�Uu_��Q>KIM�8K��bߕ=d4�>�P�=P�=�9�<�1=���=��+�2���v��t�>,Y�=1씽�H���{�7�׽�E�����⊾�>>`�4>e=>���;�æ<���=�ٔ���U�Q>{}J�W����l >� =Mڷ=a>�J�2��>��� ��9�R��7F��2x��@�=%��>�䪽������� ۾@�>�Qj>FK��72>��=-��=�r�=t��tP�>�"=D½��2�jKE>���<ˏ�s�%>󨠽�/>��)���˼|�=�%Ӿg�V�����t>�CF>�ă>ܬ>������=>�V=�0^>%v������E��=�e�56m>]�=.�=�Ԇ�Y�>j�[>�'��\D`>�o�\��X;n=�&�s
(�W �tS=��Æ�2��߹ϼ��;�-��=�eC���/�qU<	�����f����>8?�>� བ�~=�:�=��>�DC�m�'���ҾA�=&�����=D����Ľڊ==#��<'���J���E���W�>���[���}OB>�7>�Ѩ�Ḓ�U�=�{��Y���"V=z(>��1�l���k%�>�����~���5�>�*�=w6v�����?=$��=s�= �u�o��FL�=gګ=pcM>d��D����.=�Xe>H��>Z��=���=B�>>[���,m]={�j>�6>X�>-��<�>)���/�׮b>�<��>R��&t�MV��r�C=��U��Eɽ�<>�x>Y{�=�87����s��͊r�.�=W����w�=����/Jd��y�=�5���%���>��y=;q.=d,=�@U�=��=9V��85�>;�}O���2�=	�q'���c,=�t=ț��n��=�엾�l�<z�.���[>3ĳ;����	��;D8>���=&
�>�t>q�Y�p��a�=�"�>'"�<~Yc����=�P>�м,�����<����נ�=R��,��-k=�Ó<>��j�h��<ķ>O O��B4>"י�&�I���r��n��Ӗ=���m"�G"g>� ��=�
������н�AG>	��
>u刽��ͽqV�=CD�=#O���ܻ|�=> ��a�;*�=�Bܼ��ҽZ-�=/Zt=�h?ut�>�[�JZ�=�y�=�/>�=_*R>?��>?Xo>��>=eѼZ�0iu��[$=������摽GW�<�f�=��=��B>�q=/�>5T��L���6H#>�ҫ��b>��=�.�*��=F[�>������Tz� M��)k:�:���WѼn���j�>W��=�U���敾B^Q>�ds>���z<3s���L���>>}s��^yͼ��$>��������-�;k�>S��[�`���L��v�t^F�*9=?�g>Z�_>�k`>xK�>�ʖ>�B�>�t��fP7>]Sh<��u>CF<������=&;���=s��=Jd2=�s���<=��&�R
��-������)�=rv��w�7�:�5�>f�J=�wŽ,'�]9^>��g��_>�N>[���Ľy�\��#=�K=l6ܽ0xB>�J��7>!q�>-���Ȯ�>[�>�n;=�$J>�Ǻ=���1t��Z����=�b?�{#��7�=�鳹�!�=`��=�3>�A��+�1�
�?��'���z侄	5>�[>�M����2;�ҽ�`6��`ջ��>�Pw<��ɽ5S�<���bw#>��L>q>���R�J=��!=�>`4�����%���>�~�;JH�=Y��<#�==�,��WO>/ "�p=��#���0>�	�� �=T��=� >]3�>nO'�N@�>>�)��5���Z�O��;�>ܭ��3�>X����� <��)��d�>ww%�3Y�=��<����=�:�=���e�Ke>;�; J>��6>
Q���J��#B>G#ξ��C���L>��d�zL���8��龾�̯;��潳�Q�sҽ�'�.�l����i��r���\���0�6p�7��y���me>'�Ⱦ�z̽/
�<����K/\�n�$=���=>l��ʛ�*�a�.��=�q�>�(;9�(>KS���˽���&�=ܥj�2¾ ��>Xt˼�f�<~�#�u��=n�=��2���<a�����=�lb<��Ȼ>�.��N����=�k��G�>�>�j��YW�r˷=ؤ�=���=;�'>,Ŋ>�G˽�����}��c>J�r��5���`=@������2y�_(U>b��>f���A��i��<���Or�T�%�0����6�=�Pżh,4>���x�=:��=i�=t�;>��<>��"=��=@J�=�K�=�X>t�9><H>>=j����>U��������P�>r�Y=d`�=��B=�NN=�w�~�N��R�����xԄ:����ឬ�ҹ=1�a=XwC�;<o>!D=Aꂽ_�����C>���=w��=&\0�v|�<�M��=���Y��zm�vA�=I�ڽ+a>��6=���+�1�F�l+��*=���Ѿ��b=��>��0>�(&>X��R=u?j>��=�p��F>��+>�ƽh4��\d>��3�+���6���=�>s� >�̀>_d5>�α=�y�=Q�{=����9��S�-�Q^�=��i� ��=پ伒;Tt=S�>P~�~v�#5 ��A'��֛>DmI>�~�=k��ὖ�>�r�>"����]>������ؾ�؊=;�ν�b���x+>��c>�W>@��}0_=}�q>���D߼�O�=τU��-�>�&>�ǩ������/ܽp'��o?��Fo>���=�഼vU�s8j��:�>0=>�����;5����=O��P �����B[>0S'>^&N�i9��!��=7���^�=I=�C�	��z<�Yn�=�X�g���=Z�#>���>2����Cu�ϰ�>���(�\>D˂>g��=wF�=�mC����>?�ټЁ����P>5�=Š%=��>ͧw;ө>/b�����6�<�~׽�z
>�N��w�����=�`�=�#A>�s�=�ݔ�ԝ>�>��"�Y��>���=|��DN�>�-��΁>w���=�y)>��ļ4٠�\�=٪׼��[�CRнz�#>ZV�<T��<����n���/�̽����'�>��m����>�ڽ����ƽ"ą�>ݓ���9>�>D�=���>*B=���=��:>D�>W4|�-�{>6,��.�=��>����N����_���<>�-�>�@%<��)>e/>>�<��6<UQ�� K�>�1�!�@>�#��W]�>Q?d=��l5=T-	>�F�2��=�浾�l�<��$<	Q >A&����z��9>��>N�J��m�����=4��(�;?��=]����s>@w=$M,�R�+��˼#D>�ߡ=5)�=���=h_C>��� 3����=�j�5+�=�0��
�4�.pX>S�!?s>h%��������N��=����0�=:��>Z�{=�/*=e�����y=۝�_�7=��-��=r�|Z�>$G�G�>S=O�����;>^�>�v���K����Y���=>T7�>�i>N�t��+�<�6=��B>L�=�����-��Ԝ=��#�\���4��=,"�=�b�~�>?�d>�z>'	��^n�e#l�ҰM�^_���>-c=`D��}+�,�L����/�o�=�e`�P��>�-��1�=��>��`V�>���S�=��=>,β��pz>~+8��%>C`�������=��>��A�T'E�|M��|�=�x�=%�>�k}>�e�=���W��=�]���}�k��>ÇE�G�>���=ͤ$��c)=ǽM���|=L���0�>7)<�<��������<�$U=<P��C<�c��=�%]=�9�<����4f=s�=�T,�F�����6�:�>�*�=�*�>�V1����(!�%u�(jE>�8j�4�#>N>R �={�۽k�>�>U�#>���0�$<G�;��u���Щ>����"�=����Z�5>?o��	%=��)�ȟ=��=��)>��z��6�6')=0O=��㽕v�pɛ��˔>|�(>1�b=?/�=�.L=܄a>�I<@뾂�ֽ���2l���t>Z$�=j���U1�=�Ͻh7���?>�^��Z�ھ����X$�!���1M>�j��M(��j>���=�4�>╝�����X����JC��2>�u��D=��Hܺ�~�=a��;7�z���K=kW$���=���>���=҅��{ƽ��m>�#=3�$>��ν�_ɽ׀=�5�=1I�>�K=>2n��.>O}��r��<ٽI	A��{�=��ޢ�>@+�����z�4=	��>Ӗ�A���v�;be�=:�3>Z�˽���>Tn"����<�W����
�����㊾=R*>!��=���<8�=��f�#��>��>�'5�"4�>��l)�>-�\�����xZ�=��q��9�<h�'�8��<��c���Q>P�Ľ�B)=b�>p�=t�'��^C�?֥=��罻��<�
ؽ��= �����9Wo>�V=y��=\�/>[�">F�����<):C=��b=�9��g�>`v]���>�(#>�7�>��>6��>��3>[��=eEA>���>�(��4��D%�m�1>�Ǭ=�ȭ=�+彸���P�>Q]���K���꽕I!<9q`�r/�<�gO��� �nGG�Lݽ�(�> �ӽ4��g>Wl>�&�/��x���k��B��D
>a��=i9>*���S9�"�P=P����̽%&�	*u�,�Z>j��o�ֽ4ӏ�o��=�Z�d�#>��ɾ��k<e�>�.>A���Z�o<>dB�����l��=}fO>,]�>W�s��6R�����`����=�"a��B�����ru>&O���Ĩ=|B>�EȽ,�>�ۆ>֩��G��-=V}1>ɜὮ5����B>��=���õ������,��c�>��$Q���]]�\��=���>i�>���Z	�=[H�>C$y����<"��<"B<�&�=_D�=�"ݽ�@ؾ��<r�&i��7��<J{7�=�v�>��>��^=�7@>tV��3�>i��=�Q��{L�c���$ʥ��&�=v������3�t�3�C>'>Xr!>�0>p�>�X�=��Ⱦ�E���F>E��=����.I>D�,�\.�mg�D������=��>56o=�<н��~�E�-> �[R���e���`<���;�G>d�Ͻ�����W>��J�շ�=�g�>��g��|>|�> >�)E=:({>�y����� �!޵=p��=�\�=x��=���ʪ7>�-p>�SD=$Db�K�|>V�\<E�=�v<����P=yr�J`(>����L��>i�F>/�h�ZC��0>����j>���+���L�+OϽ�"�=r^�=��b��Xs=i_�=`�����=�(�>�I��8��X�>�r$�ǻf�/��d=���4g<�ѷ=Q@N����
㩽�2s>'^�L���6��0�n�e�&>�h;���>�h���>(RA<�6>8l\=ac>�%��Ek��Ð*���=y�<��D���>8�ν���>�>6h�<݈�>7!��a���/�Y惼�^���T-�vg�=�J/�:���Yi>[��<����jJw>�&4>33e����=>s&�t���¸��ؾ���=�xl= e}���o�ze�==- ��>M�>��n���=>��=ܝ<�3X�>��R��0�>`�Ƚ��@��-�<�P��C����S�B��<0�<�l_=Z�_=`W�=�&>���=΢_�Nl��w4��Ŝ�>��=������>���>�&q��m>��ӽ>>��Ӿ�!-���=W���jG>�g/=���=��=�wT=fK>�r=t��@�<�|�;���=,4s>ϩ{�xX=ڰ���=�<�,I<�%>:ՙ=>*�=Pt ���ǽ�P�=Y�S=�� >ť5��'�>�:^������%�*�r>��j=,���Բ9���=�YC�`d>/Z���/��2}�>������R��=���=��=�Ӟ>� ܽـ1=�r��u�=^C�ފ���^�C4��Ú�>�����qғ�Xݐ>����>1a<�=�=�콉$�FѼ�,�<�4�;	Fw=h)�q}q(hhh(KK KKtqhh	h
hh�ub7]����3 �H��Xp7������ ���7�Ӡ7>��������'�[}����28w���D�r�}�o7y©68����/8�ȷJ�"��\�6���Pmd��7�ε�\%�_v,��7)��C+2MX7h)�q}q(hhh(KKK K@tqhh	h
hh�ub�#{>S�W���=j��=W4����];l/�=�ټ�惽G�m>��=�S;>}��=3(���e��[=���=�\��!ڄ�ĵ�U*���ڽ����T׼��=oN>�
��NE����8>�G=�sU�d���:���[��qA����=/�=����<󃊾S/=�{�<dAۻ�E�!5J��l=�����'�=�'�B�=d�ͻ�;O=6'G>��	�>��>�9>U��=���K�4=�$�'U=k���c:�<Fs��(�>F��F7�=F� >�����#���1�/��7=�6���%9�=���f�v�\�ǽV5�=_�R>V��>���>���xl�����=Տ�<x�>2/�= ��=	�>-���>��=X�X�>p>�T����@�l�{>������+=C�T�ꪊ�8�y�w���0j��e>՛	���k� Խ��;�"ʗ�{�3>2�Z=�^��wky>��b>nѪ=��ỄM<I��`J�==K=��<UI�>��o�x�R��(k���Z8==Α��!�>� r=�x�?2�=�[!�|�5>Q�$<S��<�;��u>X�H���R=?SA��v�EN>&��=�=�>�R�<��=�Lz<W�3=��=���=���v�>�*>r��J��6L>Co�B�9<�=��&�G�oJ�C�G��i*<8>��ɹ�%�={�>>�m����{>Pη=�t���н�ɽ��=sX�� ������=�y�<4k�<E���vi=A?/��z0�B5H>O謼--A>��=?�}=�o����09Ž X���-�=�b��|{���Y=Me�<���<��#>/�����5]����=p��=F�;yg\<�v�=�j�=�E��5_f>�Y>�}A�l�)����>k��lO��z=;�>��R>� ����=8C�=9��=�ԇ�)��&)����>�K���;>�O����G<7	���5���#�$8�X�j��Q>N�P�[>B>�a��w�)<P�=r��=4����;nk��x���~�2>����c�=�]��u���<��>9=:���n�Ŗ4=Y��:�4��ex�[X�E����Tһ\
>�`>r8�<�/���`��R/>c�,�]�h��>D���2;�O>c���;�=(�=>�A>Q!Ƚu0���=v��8�m�*�)���J=CRn>w�=>E�'���?���>�pU�<1�=��=��>���>͗���d�=qA>�
>h`|=���=�E$���d�{䆼,
V=~+> �����;�N>�����^	����<�
=̼:�)������
�>�ݮ�j��=	/=��#�LhY��G���z�1gi��Ow��ֺ��i���A����G=np
�TBG�$��s4��a����t]�=\5�� )�j��=���6(=��ڽ���=���=�GT���z�ڄ9�\t��2�}�!=,�<�����<;�=�y�;6�W;ahh���1�3R=PB?=/U����;+�>G)�<�$ֽ�n~=y��yj�)�=0F#=�S۽���?j�=�>l���~��=��=��#�c�=���.��q�R���>h<�N�x�wI�A:*�,��;ͦ�=����"�=�5>��<O2����=�=����_>*��wv>j=5�=��e<�8U�*x�=s��=cQ>w��=������o��>D�=m=xA?��&�>��I�;>-�	ń�b�\=Ӯ�<����E;��B�i0�`m8�s�=V��=G���6�=H���F�=�Cf��D�< Y�<�D�>���`ڄ>��=��
�?y��3^��<迠�ϱ=�fr��~�=�ཪ����H >z�g��3彅-x���=�d���o��@�����=�<�n�>����O)��0z�"��$��=0�=\t=<�O�V��9#��˯={�>�_8�1�<�嫽a7����m7t����>���=~%<�7Y=���=�k;=��; �-=\����=T�>2ҽ!�̽�c>��5=��*>��G�ipսC�N��]��)�=��&��Fd>�۹=B�ݼ�=�  ��	�=��������	�<���:�k�<�v�=i��}�L>�>
j�Ha5=F3�=.�=̇�;��<x3��WZ=ZO�<��F>T��㌂���>��+>)��=3I[<rk�<��=��$=��>��A��YU�3`�;������/��0��H:���>y�޽e�^&>> ��ɼm=L��#��,�D�hWy��1���1<�Q>� �=�)��J�>A�J>$%ƽ��>�En<0��=N�=ǑD��U>K��8��!T>!B����>�\����Ca�=�B�=��½��?<"^��v�� \=C��\pżƽ"O�=.�=��ֽe����]=*���ݼ�n�F3w�/���\	x=T΄=�*�<+h���*>D鸽��=��=1�ȼἻ//<���=7�������;o>�>>͆/<濟=F}=��Z�q=E>��߉�-�;&�~>��>�;����5�n�!=:�Q>>�� 8l:�c�=O�"=��e����=X������=j�x�8��=�;=�8�+>�;TOb=V+�W\I=\������?=�G-���b=��B�~> >��Q��V���F<��=4����G��Q��=�>f
�=>^=�"?�FӤ<�E:�G=;�%�=|F�=���=B�m�S�<��z�;A�����>>ۍ���>/�
=�.3>����ʭ�>H��ތ.�sD�r�>q��=R0��h>He�>��<�:=A{�<A�@��a���A���V�=�Ѱ=�7�=Ȼ-�X�=s? ���޽H">�L�=|���l�<��V>#-<%h�<�=�����d>�K|��Q� �=p(�������=-�>��w>�|E;!g��1[߼f�>?��=��w>n��;<x>鯘>�T�ЬO=�^��C��!����x=<K��7�����1=ަ���<�7>8���KW���\>����<�=[>sW+=�Uj��R*�y�=p��2WV���=�����<}��=�|�D�=�OR��F�m��%�z>��N���<�#��m0=鈉�ˆ	�K�.>�ʼ��=�����Y=#>7iֽ���<��ϽUD����=>�>o@=u��=��Z>6>8��=el�j����}���oP=%�R>,f9����3�{:�%>�Hd�$=4p��+�>X�^��@V>��>�i>2��=%&=6X>�,��v�<���\！���dt>ozp���>Z�G� �'�c��=�c�<�A��4�>f���<�;�=c�Ļ?�E>��D�q
�=k�=�G����=7D�=+�-�M����f��I��� �=I�=.�C>�����h9��->�q>�g>q>J�>5�=cb�=3��=��=Fy�=4�k��ٽ+�b=��(��x
=ƻ�����%�݃+�'����h;Ӂ�����|�=���t������=�)��s�>���[�=뻽B���p�<7�p=���=_��E<;��-��>W>¾d=Nl���y�U�>M[2�jݻ����>�o�=󪰽U~.<Wź=�3����53�=>BИ�tņ=���=$Q>�3u��<�J�����=�c��jνSޛ��Xֽ:�i�9�=�!:>��;>[�
���>.Ž�]��Ӷ������v>͎�=:=V=}6����������RX����4�4���C=_����@k<ꡬ��=R=�Ӟ<3���<*l=�&> ��=z7*�Mۢ=�T��J��tb�<����G�v�&�`�}=��T=.>���$�7>i�+���|�I�=��2��S	>�h>��}�4��=&��2�Y�YJ�>I�E=S߉��c½0�1<�_�<g턾@�`�c� �R@���c���dŏ���,��=ې/��9�<j^���s;�Fx�w�&�7,0=�N�>���=P��J"Žz�R>�Л��>Y3>�
�=r��	+���!���ϩ�0�0=���>�7������<�Y���� =���=տ��t,>��=�#�H S>s�=�!>�]A���ʽ��/>'D��+��c�<�o��� =�p���6y=�5;����=��۽�S}����A���C���	��.v>}<t>c	^���i>�9�=�
3������z�����=���X��J[U>"f����7>U��=�"�����6�=�k�=��=s��@6ڽ��<�= �<��_=��=t��`��=�G@>`?�=	z= @>��;�LԽ���2u>Q�=��[=Y�4�Ќe=�[�]����W]��ׁ�rj[��B�AD�=e	>$N#>��>����xn��^?<Ƌ�< s������]�������$�=`a��Hz�M����9ν��ݼ z�=�K��\�=��`>��B�y�=�^�
<��<�N>�h�<�'����>E>>�<Zϧ����=?򛽟fL�`�:�py>,V=��$>�yI�Ο��Q�>�0�=���mᇽ��#<�&��i�=��%��j=�&%>�7;�x��woG�� h�i���I����=�ƥ����<`�1>�.=#����N�=L=���e�=ީ�=���<Ll��e����<'�־��;�F\��q��=y>K�=�FK�1�%=�E<�j�=��<:]1�2½��-� .<���=I����=ŧ</�<�ޑ>P6�=�<���;퓰��e�5��=9�=&w罺�>���8�=H��g��<	��=&��<������=,N�=p�˽��[�2Y�>�e���� ݢ=���=ZL�>��佢����m>/�>;��&��>�_��d���}�N =$��ם��b�=T�k���=����>��=i��1ʖ��ܤ���Ƽ[?��c�<��d=Ç=/�M>�d=>��y`8��v��/��t�6���b>Ek��|���	?���=(��=����r=&;���f=�r��ϼ4B��Q;"���==�^7=��%�xyȾo>ܙR������=	3>z�M�c=ṽ��)����=.�<��@>�>��(_����Q��n�5/�c�S=����c����w��!���>�=v�����=��:;Nkw�K�=�z:>�?�=c1�r��;���}=���=�@=�I����8>��^�s�S;�0>T�D�M�=pɾ̜�=�1>i������=��I=_[�2m���g?=�s��>X�>�z&>[&�����<! ���5�{@�W����=�E��Ip>N|���=l6k�G_!>��˽R�=8U8�B����>����QY���`>�䒼D�c�b6F�s̍�ȟ���὘l�l��=/�:���������� F=�B�����=1>tє;5T=&��<
��W;����:�V>�%I>�D�<�󿺉.K�����~͓>�.?�+R=kk�=��'=�D�=Mܼ�A{=��=�->[*L��7>݈�<����t[>����"z�=l��3��<��(>q)���=���j�;�
�_�>�>�>��_>{=W��=�φ>�=�	)���=؆I=�E����<C�G��h��l�=_�>��̽��彂&+>�"��,��=�s�;8G>"\&���3�^?��;Q=��'>�y���#=�^���d>,�=b~{��/���}F�=l�>��<e��
ͫ�Q\*�D�<LM=�=eRL>�[U�1*(�Ͳ<>�咽g�=���i��\��I��+%��+)*;;lK���n>�	�=P���/j�O�<n�7������3�稱���>�J=N�
=NE=��!�G��T;��m>��>8>�;�;�ݽ�q����=х�@@+=�b<��?�����@��㏽�=�<�H����;����/�7\ =��T[�<#n�����=g���%u⺛(�=F��<�ϡ=�m.��N��8\>��#<�R���L>vKi�S�c�o�T>�k��(5>_�+<=m��bT���J �N�>ϷO>(%Y�j���D��=8!ʽI�=b�޼�9��k�C>&>�Ѹ�B>�S#�����H=Xo�<Ec=���<Cd�<��>4�>���}Y�>���=m�w���9>؏�S�=���=E�������w
={=*N�=y�˽n��������>��ؽ��:�!^=f3_�[��c�=^F�u>��1>��<��>�Φ=�i��~{����j<*�<D�3�F7?�·�=-Ǆ==}#>� ��6����<>��<،=�B�="
1=�
�=�~<�6�Љ<��ݽ
�ּ@A=���=)>ɗC>40���T��(���p�Gi��� �=��żM(���z:o�����<A`>��>:�:)[�]
}<��+<�7�.�����KN-�����愽�d>ق >��(>�Uj=��>�V�=����_
�g$�� 0�x�:��=���G��ˠ=v1��]���f�=AB>?V>>��E��M�%=��=�u���G�J$��b�>6�� ���.=8=m9�oP=�R��T	>qȷ��i>���=;:Ƽ�T	<er@>-�=p���`ú=D�\�CQ����;�/��"����=��>�.��l�=�g�>�JW=���<�6>mW�=nN �e��V�c=~J�<�O&�4�۽�2�>��D�Hp�r"���zR>=V�=%4���q������g=��h<lx=�ޯ=����*��=���=�P>]n=-Kٽ�,M>U��=��y�m�I=dG>�f�<9��=}��>7����ֽ��=�~� �3>	[�=���=�۟=+1 ������9�=#��E"">?6ս��.>�M���-����d��C����y!<ĝ����q���a=e,�*K���>k����pk��Rd>�ɫ�(���(Y>r!����&I���7<G3�s��=����T�e�>Vs�A�=��m>L%ý�^�<[���)<�8��^݌=S��x\�=C���ё�T��0�b>�<�<%L�����Io�lg/:�)b<�\�=��=���q>93�=k_�Y��&�����J�=i9a>���3[*=U�=��A�tc�>��9��<v��_k=�[T=����׊����m��)���>3[��|�<GL=�p�=!�f�2��=@���0��fa�>uΗ:�v��`=��d=��3>Y�l>͎=�Ž<��t1=��=�˓=�l��;	�u'���U�=�j> �#=���=��=R�y�o���}���P��=zD����~�����Y9�ԁ�=��λ��	�`齼���*���l�_.ݺ#��>Q�#����=��=��D;�c��r��7ǽ���=:N�>=���m�=��e��a�� ]>F��>M��}��Rl\>��=��=��0;[�i=�A�<I�<U�Ž�7�=�@��#a<��� �`z���PO>2ϗ��/ݽ]@_�/v�<�>|��=�U�"��=R}�����<�v�5:�<�1��}�>Y�
>�<��l�b!���>�o�6���F���n�=�楽b��Z</��=�W��n���ɽÈ>��>b�Y>��5�δ�=H�Q�%M <#hż?��g������=�`�=�R�,���^=j�I>���=	b�=?��E8->`�ٽk$ǽ	��^d���&?>��@=��U<=����m�=�y_>�����X�C������<tJ/<�(�=aݜ=�>'*V���a>6k���P�9��{<d�3>��U�MQv=����� �S>͹N>�ߖ:&��=�	=v�(=��6�FƗ���߼�DĽ���=��B> �m��5���f��j����Z0>�ç�NI�=�>�iG��=P=�нc�=X���9�S>i$/��{�=�6>y�J�Q>ϙ=��;>¹E��Q�<|���R�����X����C��m<�v=L�½|+�>���={ї>}�.>��<�h߽;���va�3�Q���:�|F������ҽa�S����:��;_���7�=�T�>-���5��;c����F>x�T���(��=�f�=���U6��	A��A������a�v��=�ۺ�1YϽH\���L�5f�P�*��A�=�x�=N�0=� �=�p�>Qzd�r3�=ǅ�<*����]���u�wd�=�P4=�:���3����ϻ?3U���x��$c�)�U=���p��ϫ;�wTo��S�=	�w>�%k���9��i��!;>��>�Yb�;��=�3�=*=���+>R@>�%2�H�u={���,�=SXj�2�-�K����0���H�״�=	s��hS(>���=F��>���(\\�d��=+�a��%����C>�O�=>���>� <��/=�B&�e�=���<w�<�o�1�q�+�Z>$h�}h&�잣�Qhڽ�����1>��=Ɋ3�}��Zm/=�a���	�}�½J8��y�0>�^n=kE>�EU�iE��������n=��a��34>S�->"��=Y�V�D����9=++>:�<D�W>?�<Hnսs�y>��=��$=�Z�j�!=|�/��_t�DѼ.y����=K�ٽ/��\z�=fb��P��EJ<Ð�=W�?>3�S<Q��=c����
��_�<������==�>Z> ��� ��D0�=p��=��h�&=Cu>�ν8��=�X��U󿼕A�=v�=�:9=8:"�7������s
���=�9<�����i��!��=�8y��(=<�P>7����&��0>N��pGN>%&��L$�l�����=d�Z��U'>`�*>��k=����}�=��,��9�<��>��8���=]�=q�<{���r?�G�"=�mR=�f�>��ڼBϯ��Cn�]I�=C7��_�=�s��,ȡ�����sv��/��);#�>���=��>FV.�����f�E>�t�>Q�W=2x`���<=�9=��P=��8>�σ�
2��=�;��:\�J�D�r� ��1�<��=G翺�Ғ>=�ȹ7,>�=�F���,�2=]=�=�Q>�nϽ�C���#>��>u�/=^;�=�y༉��]:>��U=�D�<ăU>��%=^��t!>u<�wd���꽂\���T��g�jpH���սg
�=�`�a`;��=%�`��3==�5>u�{>��>��B=s7;M��=ߧ>�h�>������=O�5>�ڼ<�^�<��=��u�u��YC��½���b��=v`6>�!�}��<X�>��K���ֽ��>>�x+=G��=��a��7��v;��P�ƽ<�=spY=�Į=d0S>X���J�
��������=/V{>7S�>����N��<�	F��ո��E�=����/�=��*�!��<?�&���>����X��D>����-���Z�X�
=#Y�=�S�z���B&���~=�8�<ń4>�[����O>θ��0������������BF���L=�bC>ؼ0�H�WXD=��=����lU��aE�;� ���:���~�>�>�=����=U5�<s��=�v�=�	t:6ݺ=��M;�h�ʁ><N��PK�Mh��(7��A�!���J콣X�=���=�S��yZ�=�c=�M���=��:<�=��Y� 49>�?a=z��=�j>��=X� a>�o�>
��=��U�����8P=��w�[ԯ;�jQ�ip����;)���.w>�-"�������=-k�9T�R��E��}�gf�<�9��ɏ�o�u���>F���k.�w�K�U���o=�9�=d�<ף׼XY>!��B�>��>a�4>F���}>>��@>z]�����=@l�!��<�s����<{7��_�=J�>v��)�=�κ=��=�<�|�e=~���D�=<�<9�y=�k�����<��j���w�x�=�>���EB3>���<�E���2<����R>m��;��=�	=dǑ=z��=��*=�"z��$��Ҙ�=U�C>�]׽�=���X��T�=�wY<�������h�=^{�=7C>�沽�Ƭ�l�Q�">�ݼC�W���/>0OF��j�x�Z�X!3<"E� �>�>>�`�=}��G�=8 ҼYe�<��N�+;�>�	�=S�B�(�iC��U�����ܼE��>����$V����4>X��@��࣍�J<U����=%�=?� (<-����Y>su��&��T�ܘr�D��=8>¾)�g����N�O�\��T`=k:4�-j�X�7>�3=7�.=T>�v->�Z�<��>��a��-�z��!='�����>׸�<5K"���^���>�$k���SE)>w�}=|�=��s<\���>�g1�N�Ƚ�,��g&=�e�@���pL�=e�����K����<�w}>��z�]a���O��.�x�'Wѽ_�$����;5ȼ=�U����l�>��>0h=G��E�>>X��-2=y�K�O%ܽ�$���Q<��%�x�ŽmC���՞�
1�I�w����=�("=�N�;�5;>f��=�����=W/�o'���<9�.�!-ǽn닽�����˽Ԇ�=a�����-����=(��<av2��g=�0>B=�l�=�Y�mL��d!M>�T	>����Ŝ4<Y�>�,I���Ľ�����=���E�-���=��;=ZS��+�hw���x���K=y�+<��<�e�4���/�h=�����?=�_}���'�U�=�=��q\�=A�#����+L�<ףi����֮^��CԾ�E�;q#=i?̻Sg�>a���||�����/;�ǽB׽�r>����jX<�ӭ�t*��]��?!>�������&J�=!��<!�(�L�J�n{��Ю�0���ٚ1<?1߽�E�%�����͢V�������m>R�> ��;5
<۾x>��N����=�/;&�C�����Q���粺=��ؼ5�[�4ZO���ü���Դ��=�<��=�>ڄ �/�>�Ƙ�[>�
�:9>�����{';h{!��,;>�ֽ{k���V��2�7���;����<�)O<2����.{���=L��<'|�_�I>��~;����Ž]+ҽ��=���.�o>�A���=������S=�D�=A�= ��=I�	�%��;=]#=��=��=��껃Kd�Px�<�
N>�X
�l�l=b�*=�-�<D�7�)~7=��W�k-F�I�=�|���o=1�0>%��=�W��E����#>̖���=��H=��0��pW>d-�]���Ҍ!<7�+���=G˽4�Jf�=��[�����>󱲽�#��T"=X ��->6�z�=��
>}\���8=��=��,�����_�=dk����h��Ҋ=8줾��=�D��N=�=�����>��7��������`5�=�}o�V帾ȫ�5o���=�^�=�Í�r�=�S<�=���= �I��n>
�����u�=�;=��>�F5>�7-��mt��-���7>���x�+=���=!.����e<[��9�X�\�=A�z=u�C>�P@�qS�=]*����x6��F>�[�|�Z���Q����k$�n�l��0�<"���T�>�_"��0�=c�k�㠻�XD����<!�=�>�CI>��<�.�=��>�=6>�,�����=9��<LY���f<F�<�6���=�f>�*��uE=x;�F�����N�:=�}��3 =�g�=	�>]!=�%#>�k+>W�L=��3>��ɽ�[=���ֽ7�l��>�&��U�}= �>6��;0��>���E�=b�H=>x�<{O[����=�r=�)���Ow"��rּ�C��E�<��D> [=�3�y*�<^V�ri-�"�<D�>P|���^��y�����Yps�&���1���|>%n,>�F���=��>े=3��ˊ\���ڽ�Ͻ�-e=�H�=�E>�@�<��?Fs�Nw>`�\�t?/�>*�A�	%+>����4�j>��
��u���Oe�ħ>��=}B��)-M�n��=V��a��=@�Q�_:b���J�2gb=���=���=��<oGc���>�B��g�>�w*����{����=v����� Rн��=��=�aw�,�i������=�fŀ>��c�.ww<�]ͽ�[�eԲ<�H�;X|z��ʁ=Fv���
��Bq�����'��#*����SQ��u>�]=6F�[�˽�靽��,�w�>��X=�R���Ľ�*1;y�6�o>�;s�G�a=���=�R�='Z۽"vM<=��F�> ��=��=m2~=@�:>�U9>KP*��0��*�� *�=�ʋ>��>>�6��s��9@�%>����tgۻ��X=Y�=�ˍ���(�e�~=]��=�r=sy�z��=�{#��D���3��"��y1=�Yн�P�=nTJ��0���|���<[�B���'=^�μ�e���l=(�-= �->K��=5�>���<#\*>=k�=�=�vtq<�Ľ��'>��
>�ҽ�~>�����O����>�����<=n�>إҽ)*g=BM=x�;�S�<h>6.��q,�!��Yh�<�>=��<��_WۼU�R>>��>���*�=O���z� :�=\�4밽6�eNm>�j���hսV_>Ry����=�ʺ؈��9�H�~>�:�<y$�=�O����>E�>���7�U7�<��=w�4�Gf�o��=~��=OF3=��@��t�7�>>�	�<Ө(��۽�n�����������\&D=
�=��½A	>��>r��<7���ʮ��x �ƛm=�>��[= *��4�=jډ=�$��B�=�����3��e�=3_�r X>#0�wο�����?�R;	<�=�2;�J�=�r�<X������&_4�O��=x՗�r==�=�=7)Y>n�?�)�M��>>���C/6>.���C<�ǁ=؉ļ�K�=���B�>���<5R�>���=k��7�WX<C&�=X 
>Cv��/'.>g?i����m*=�Y�=�
�8��=�K�=��=��=�@��{��i½��<qc���=X��<
FV�� ]��=�	��,<��0�Zc���꽽1��&>(�8>�P�׵:�K><���X=3o�=[�=�r�
;�r�=K���2=}�>�>��Ƽ6-�?4�}�<��P=Te�=ጣ=��ǽ�mȽ�����=N򲽏 L<�YA�+�{=�@<qF��E>����򯾓�@>�}�=���=���#>4��?1�S�c�k�<J�>P=�=�4�=>��>���;��=�"�<,h>|�>>���2�J/>I=>e� ��V>ĝ�p�l�\{�=�<���<���ʷN�g�b��_��S�<��@>6cc<���=]�ӽ�>�=Z~�ͣ�=�s���=d�>�S�<"��}T6;u]�G>�����H�=�푽����x�i���E�4��Ņ�!m>x)�>-)�<��<\
��_>���O�۽�yA=��� ά�٭�l�پs�����=
��4桽�u6�W&�>E깽�5�<E �=��O=
E>�5��2�$�Y��a�!��C>9w�`�$�Z珽����g>i�=�\L�y��J/>#�)>/Z�����O >��ּn^�b�����=�ع�KW�5!"�+===oy�<�A�=>۬=�|<:�����׽�����=[��0QB����i�����>#�����=�U�>��=׭y�w��<��ܽ(��<B�ĽVl��e>�O��Z똽mX�=�ս�1X>(i3���>*M��I꽌��=iZ����=^�i�2�~b>iC�A�>���=3��=&�&�@M=<��=��(�8>(�~��l<T�>b.�=	��=Ȯ�<v���D����ԼY��<k<!>�>��fM=�BP�;��	�ܽ���=����y
>���;����ly���=���31>�l/�O�m��^
>o�[��h �����n����Y�;����.�-�N�&��'����ԕ>���=y�����c�=H^��T�=�%���д��/$���=��k>1ƥ��_�����=�.ۼ�ε=�>�=�ذ=J� =%tٽ>�P�#��=�W�=�G�t�;�Ch>T>'W�Y�7���;�>ͽu7����<5�$��BM>:� ���=@� >�ＸI �`�(�>c߽p�����7����� �*c�=���6νۨT>~ߖ�U6����(�=F�>�-��8何t@>O�ؽ��?=�߼�n�=��<�y���m�=���>�V�#�<���=��t=�����1>�z��.P<���=}Y�m�ջ5� �-t� ��	�0=SB�=a� =�l�=�g<�,>�[=�N�<2�z��?Hm��
�i��; >�H�=���*/�RE�>̝b��}
���H>�Ɂ�p�=��=�PƼ�½r���W�=�ֶ=�ѽ�Ө<.���U�=Z�D>;�u=�@=�[>z��=�d@=��=pN�����D��+Y=�ּ+%�<���Jm!�:�>>�׎=eЈ<�	*>�-)�	 ?=h?�>��X0.>6S">u�>��;�h��\�м?�<[`)<SO�=lҠ=k�>���.��n�-��e�=�{F>:	F>�i^>�8�=/_h�����4qĽ���섕>Ǳ4=�`8>%C껣�b=6���o�>}�����=iG=gA�>��<�:�9Y���=�0Z=�kX>z�z=R��=��»��-�߇�%�d>7�1�m;��mz�=�#<~�V����<p�>>r��;A���!���s��Dq���&�<z�.<�[=�==��>��<��w=Q�q���`>���@����C�s`%�IPn=5'�~�O>��<>xe3�}�j>�>:�O����'��B�=�i<iD��=�8R>�S2�y�=w�=����5��*�>)`��4<v>���;P<d�<�����ɽ�K=��Խ�"�=�=t>�뵼Yc:��Q=q?g��F��x��=���=|v��"��=b>'P>(e�*�=)u���1�>��1=���>�n��^��=���r��M-���P=�;�=xj^<}�?���I>I�*>J���z�7='`��e��<q0���>�<eVY���P�(pJ�ݶ=�~">Y[b�=ų=-]>��=�>�P=<�=�C���bR>��<�w-���^���,<cۤ�#�ƽ�����<��Z��<�		�3Ɓ�c�5=�3.>�FL>�1[>���=�~��\��+�N��&�o8�=�C�<k%J��>�C�#7��ȂF��}=H�罦�>^�+�,�Z��żس���Z+=r�l��$���=�S��I�Lt����<��&��"��+{�&�3���P|�<kP�>��>�V��t��(�j �d
�=!�i>�7������^c��+�:(#�~�v�2��{�>��J;4Z���A�����=<�z�=�>A`]=��$�1�mQ|�z/�</=q�S��.��u��<�>.[<o	��n>���=�޽���<�Ef�h�R=. ͽ�P�5�&��!3��f̽��>#e��L��=���֐=��>��=4n�=��� G�*-B=��+<`�=_�6;�M:��y
>��<�'t���K>Y�w<����l}>^o#=�~>��s>HT$>����e�=�U���X8�����8�̵�=:j'=�{�=��=���=�ҽ�:��(�#>4\M=u��=�tŽ��L<u��>BƐ=De�ř�E�=�������h�<��=lký�`>LI9>w6���<D��;:���&&��A���=��ż+M�=�pW����[ln�4��"�P��݋>C�=@$>Oc�=�"�=>k���cȼ&��da8>�e,>�k=���=�7��B >(g��&��>cr�<K��/�i=Q�B���8>2	�=�>�����.R<掝=���<��3�u_,<R�=���6>j�>V]����=���=�������+'��~%>�.�9&.�h*�%1.�5!�=,��>FG�EU>���=os>B9��`=D���mJ:"I�< ӆ�t��=�G�<�/�;g�>RB'>�U1>Hש�,%�=�$N�$�=ҞH>JF�����<�_��#_�Zy ��%�k��>LA>��X>"�=&�����=G
��})O��=���}B��ȱ��jB>�B���=�-+� h[�[dZ�w�~�1C-�ȼ[=b{�=��=��B����g�>�>���>N=��U=y%>�/k=SV�=u�<���D">��6�$�=:䒽M�j� �I��!�p6=!�c=XJ9�f���.��=�R;>�H%>}�w=�=Uн���;7�-�ʔ�=؛��R;M���D�ts4�X�>EB4������<*C�T*> ~����=�9�T	���T�+��<-��?U�=�G?�k�޸{��;b�C>�����c콻Wa�@�=[
<75=c�W�QH<]��>���:-F�����4>�L_�h��{>�s�O6>��<:K=e��=�L?=U���6=�GM�\�=9`�=��Ի�D��6(�=:Z�=�=wAH>�S>Ĺ��d���ٲ��Q�=�����==翃�(詼�n½�Ͻ}�	�oF�=DL*>ܟe=q�=���=V{ý9ࢽ�w=1��������]�;����o>9��=���=��I�<��٫���Sh>|7�>���Q޽+W=q=�?+�!�`��9:;NW���@��@�^=�-��2�m=2 =����֗�C	>p�!��PO�7��<�����E3> Wؽa? <�QD>��8���>%a�<�6I=���=7^��"B�=w�����<
p<�6���w;�h�H=Mc�� "'����yT�:�=_"��[���.���>�:H?T<\vK=�z���;˽�D�Mӳ�I������=���*��=o`F=����r�>��ƽ��>S�|=���=b�����>���=&o��&`>5��=`���o4��D� h_�:����o����;�!���P>��>x,ǽ��m�& � 1=��ݽ~��`1���O�<�.��˾��Mӽ(QL���C>m��9�v����n	�<��ѽ���˿N>>�Y=��=`�c:�=���=�#���콕�Խ(	ӽ������=�Ȣ;�[=�n�i����Խ!�>���<�]O=��6>�SƼ�n�>�E��3y��c">����Ŀ��%>$U-��@�=p.=�*�=#����=T�V�df*=���v���|=B:�=S_�q,;�c��j3>p=s`���<���=�>=��ý�m�:��$��<-#>&�8�����_>���=, �=b�+�U��=�4�<6t�R�|;[�;�U�=��!>~�>�!=�Y=Q���k>$ڽwT��/k=�c��!�)����\�=�j�==Dٽ�,3������^=)���ٚ�=�#��-H���=k��=g(�_�G� >�����*�ܢ�3H>_ D=����cμ�㾼��>�p�=������g��.�<s�ؽ0�=-��=A�>׿>��o�%=e��=��$=��=v#`=1,`��g�<}q��خ��S�>���#xb��j���8>7f>���<��)���<=��`���>�ڬZ�+�E�W:��=�4�zk�'a�I�v=�J��Q�>�����zB��T4>;@">ϳ>�ȼ�6�|�<�t��>�C���M�.z&=��{��,�=�\Z��Y!�#�[>�>�	V<�A�򜽀��>\Ö������0!>-`g�<�=_W ����>��=�K=��<=�GĽ=v��e�ü�|+����L�!�Xz@����@Y��Z�k=�a�<��~� .>��1[�<N�n<)�=8��v�>�X:���=��>W,�=H����*t�= �|=�]�9=��);������^���Z�
���X<1�=|�ǽ��`��۟=����7��<�����
>),U���$��=@�=�̖=����=��=�����>7� >��.�j�J>d`#�C�\=�<��S������c��.��=����rw�>7=��P=yW�<5*>m��<��2=� �<�v�?�$>��9��t���ƽ������=��4��ٞ=�j\>AW�<	�S<�#6���� ��W���*���e���o6>����Ͻƽe�7��"���X=�>қ�<q���fq(�E�R�|43��������@�r� �<����2���j���[>�T�=2�3���?�b-V�<,����\�u����Խ�˜�a�-<N�Q=�q�=9��=Ґɽ�Tg>�p>��h�.��렄<>,=�Ő>�=�{Y�	9>n�>�B���7E>���=aH�=K,=�q����m�>�$Q=ߌP���p��u�=
l�@����=�Ͻ��>,+�=Lmټ���<��P>�~
>�X�SM��G��i���!����v���_�����W=�kg<����_���.�����=�â�=սw3Ƚ͕(�')��g�=n����O�=R^ý@��h�>�ި���+�n� �*��;�_�=�o6�{�=��]���G���>o��=�m�>aM���]�=lW+=�N��I��<��H���=�Q=�뒽�S��@�>�o�=��=�M�;w���T>�����>>f>_�V�N_=�o�ռ�9��=�S~�������?�R�;���9��>��=�ٽA$��z}Ž���;�%�=���=I�=&Լ�]�=�iԽ��>�%o�PI'>y�<x��'��<	�q>s�<2�=6��n*�x'ͽ4M�>{74���f����=Y�½��H=3�=��=��'>�tw>iIO>9�A��yY�p�>�<��u�W�,>Q�=h6��m!> ��<��� �s=-�Y>�r�<��&>��=4��;5A��vNG��=q�K�X�$dֽ�b>���=*�=��R�n䌽�Y�>��̽�Ç��ýgJ�=��= ǽ�Y=���=[��<�yZ>��伢d�=���Ғ=�UR>�0޽;�H>�ƚ;�;C��œ=�9�{��=�U��/�<Wc$��=�3���z�>�G�����<SuN���dER=�4W>��=]���W��g�<�a�=��=i����{=s��`�3��(>Ҋ��=�v�<Ж}��+<
 ���f�����vW��0��� >�߭=�">j�<gv#>��*>�w�<&�2=D����Q=�f�=۾�S1C�:$>bソ���<Ӝ(��>�F�G(9���=~�>�v��$>��B>�􎽋�<[kO>=%��:�=�V���=gC>��B��IE��g���l�=�Э���k��=���=Dʽ��,>Hj��P���s���3����=@>�p>�)�=�Au==>�y=ו>ir=�a�GN���bK�����F�>��i=��;���#Z�=3 F�9 �����4Y�=}� GC= Z��'��+Ҽ5��ʯ�!*׽��� X��_m=jZ��>?ʓ�|���I�>0�>>|[7=��w�D��6ü�Κ=a������gwҽ�b���:�����܊r����=�G�=q>ڵ�����g�=���<��D�2� =���=_��@�2�"3�o	�=�@9��R�<�K[���2<%=���=U`���C�Vb�;�װ=v@I=�M>��=�A��[)>�$=?�.�=�W���������7=#L�<�[H��;���v�`=E�U:�=߳�>�Ď�S���4�=Q�ýS-��*���<�b����h�l�r���[:W=����yB����<�y==��g���\�!_U>���;�tF��
=�}���ȁ�c��=Ur��9��=*�ͽ�'ٽ�8�>j��=��<1L�=|o�=\�U�!�v�ߔ����a�<T\�=-�!��ܶ>b��='��<�M����%e��jR
>�!彃�>�=Ka>�^L��#=H~;8����%��mռ?Y�=�!�9�>��R>��^�8_�=���L޽�_�۞F�n)�>=?
>����=
�=+Ľbh��Yr���ί=�T�;�=�LQ>ޗ��_Q>�D]�c��ڑ�������=���VUʽJB�>U�U>K>����&O��h6:>�*0��� =!�>r��$��'���c=z"����=B�=N���q�=I���N�=��b=�H�<��<>T���=)�<;7�,p�<�:@>l5��y(<u�ܽ���bH>5��>`h��*ú��>���:�=ӹ^�M����=�(��T�=�+2>��ͽ "���ѯ��ܣ� ��C:<��<���+��@��=�5�<�>�ґ=l7�=�e��'�>)'��"���=���=�E�=�а>�"#�i��\�P���H����R�p�>:�<������i
��`>FM)=��)=�r���=N >01��"�x�d>T����D�(s=>�;�=���=�2�>,�+�r�<� �>ǰ�<ƍ̻�`�Uѝ=S��<��M�맇=��+>�#9>w���t��hJ������l��	�8>&�:"=��	��^>���Z�$=�=M>W���ü��=8$�&�=���k(��bL>U�+���<�ᒽWr�<�y��be��~�=�-�C&�<��=XՖ��My�'���d���g=�۝=#��>�<k@���#�
ǂ�j�C>�J��%�~<�Q�=�6W=�:f�w�U��G�>��?=`�ҽ�@�4��<_kg��J4���=���� O��j� <�|z�����O�R<.j>|���#�:>z�<��#e<�Z.���
�Wy�%󽽤�<o�1�6(���>��0��w�=+w7>���<+E��o�=7��=lj�?;v�lQϽnJ>(J�>{�$��zX�o��=]G��-]6=��w=!b5�<s;k�N�/��=��殼�q�=ؾ���7tR=��t>:��Ps=$�Ͻbm����=�� >&\;�_Z��t�:��d>�%*>�����%>:v>��F��=�	�o��%�:�P�>[F>�߮�;�:�<�j^����%->�(�E�<%a�<4+���F!=m;�O��r�"�<��(<"��<��A��= �9>�i�=?�<��:>X t=�K�=$.��j��{'4��Xe��_�\8��y������^��;�x����<�7Ż�x�<���]&�<Ǿ�>ނ���2�B�⽀;�� ���+��=�c�<)��<�F>cv�<�����-��y>&�e>��w>�j��_�<�l=w@;�=�;jW���>~=#�<�'�=��=j9e>�m*>���>�B�=8������훼с@�N논�H�=Jt�=< ��8�S<����ǁ;`EG>�����=����t=}�W�<��>�:�A~r=b��=_U2=s���_c����>	��=AV>8��> �>��B=��P��/��5B:��M;d�>	T<ni�=��+�@=�>�=hd�=�[>#��<�>:�>ڷ��d�8]%��>��>cu"����*��N�L�'��H>��̽'� >R��<��O�=_��`���3�N�>B��=<��=)Z*�GT�>�l>�lH=��Vn��YQ��gX�8�;���=zb>�T�<C�y�����}u<EO���>Ǝ��{>���]�<���=�Լ
��=4�̻<_ٽz�
��C�����;7��=)��)���+~�>��λ)n:=�>��->���=Ŵ�=�=�=��T>~]�<6��<���=B3c=ߝs���=,Z<v\�=��T��f�=JK>i�Q=������
�c�<�G"����=>vE�#ϖ=�h���<ɐ������Vp��<^Q>|m�	�D>ʐ��� >HN<� ">Y��=�6b�<(�>�	�=9�ڻ4>�E��t�I=�|�?N�<C,���=�B>[��˗o>49p>�>:����(�%�Y�w��G��^譽ӆ$>�>�p�;�>���<�mE���^=����eL=�1:��I!>K���y_Z>	�>��c=��C�񮵽J�	��la��7E��0�>�Y>ŧ9�N�+���f=�[>}���m�>�I�aa>H�,>�i��Ԉ��f��*�B=͓=�C�=��ݽ8�;�pc=���=���=�T�=�6:\�i>�]=�x�J��==>�ȽK��=�/�h��=hi9>6j���UB��,��i�޽��=���6�%�������=��n=@E2�U��=�.��������н���=��>�3K>��=J51�o��=$e��[S��1=�3>��9�'s����'E�>&[=pZ�=��ʼ�Qܽ@F&�y��=	Κ=ouV=D�~<�>�����.�=p��j��*d��҈��C�=3'>.��>ְ;��V�r��<)�Q>�����=i����Ř9�͛v=w->��>���=M���\��]�;�G�T?ɻE�>'�˽�Yj=���=Y�L>�<yA��e�$>Y��;4qa��J���F��^s=�$=�&����(<�a<�����>u*S>�c�=0�M>෿��vf�S��o]��T��Dg>N.��V���>xon��
>�<>�#(�;*8�~�=��'�Ά����=�t^=��T=��=�0@�9.>�:��o{+=����&��{��C>=�ŝ�VP~��0U�X�=�� �$e�;� >��l��<� �
��<�>��5�6�~;@�<M�%���=���<+��=0�u���=o
���ճ=y�Z��NB�'>��j�=��r>?1Q>�/��[�U�d=k�;��y= �(����='���e�����=5M��Z�t콰�b=�*K=�,�>輡<��_�F�x�B�c�rN�=���=֑�=��Y=�Ҝ>�O��nr�<w���DԼ�����(�h�"=�zZ����=�P~=�m���#-�1�=�>�z�`u>�q�i=2��w=��i=r�:.����4�8ۜ=G�j�8N���D>��ŽX��)c%=���=#*	��>���T`>���Mۮ=���=���<T�&�[%���m��Q��V�����=Q��=��=�/��� �>6\���&�==��= ��?�<�n�Y����{=s%̽#�=㓆=Y<L����=m�<A�O���=�w0>&�=�ϵ=��+>"� �Oּ�膽��s>'f0>I+x>�Q�4��=
�>fh��"��=3��Q��=]">��~=ڃ;���=��=�(�Hç��s0��v>P��W�>=@>��Q#�=��>��V�F��*7q�S.��L�<Qe7>�f�UMU�=!��5=O�=������5������D��ՙ�����=�>̽�`>�c)�䶊���i�>!%���Z=ǎ�=>�f=�=�� ��S��e@=So����=�:�V�=bAt�ĲT=g�j�8��'L󼚏X;Z->�����9=�������I>?"V�"g���<�
��;��<F����E��3�>Z!����;1>��(x>�A�=�͐>�q==�t��p:���=���=��u�Ԫ<�&�e<��]=�=[�9��Zo�	0�>�fu�1ɋ=ܢ>���=�~��	։=_Qd><W�:��=E�=�:�=l�D=/�E��bV>�L>A@�=SkH�9�)���>#�s>�W ��>��5��/S���ֽ��)=_��=q�V>7-&�*�7�ު��k�y��=�"0=�<�=6jڽ�����Խ��'�R(����W�p"��ڬ��s�=o�Nk�ڞ�a: =0z[�	���l'�ԉf�,.�<DϪ;��	���<]WT�5�&>�>�=g�^>�]=��=��'>y�󽋃�=�R�>b�B�n.�����9aϼ���<(Џ=�C����G=��ٽ�g��y���ދ�kq����=��o�sa�$�0<#b���3K>pS>�]�=��	ؒ>�<�D=�k��'�>\><a��;���=0�=с�="��aD,�֑�=۱Y=r��ս�K����B>X�=+u���>���=}��=;u?=��Z�>�<�>ڔ�;�~�:�,Y=��?;�:���7>�l]>A���ꮽj��<���<�^Ͻ�:;>"�2>jg�N��;�`�=nu��D�3=�nP>��ܽ�o�')�=Ty��MX���=���>%w"���}J;���9�Uy0>]m6="���77=�z=F��=C�Խ�j=V��1>�=a�t���~��;�=�hz�f\%>H����*=�s�>*]�=��>4ؤ=������o=��4�컂=�J�=[g<�	=*�Ǽ���}�=�?�<�lc>���<�M.<S����x�a7�i����=sx��?b=@fԼ���=�[=���Т��2=�����>�Ժ㊲��)x޼�vQ>E%�����n!��1k<�~>˒�=g��=�ю�����E��_�������m=��=l�:�{*<L���\�=/q=�Rڼ�5�=��½�A���`����>v�V����e�=��d=i�j�v!=W��:��[>1Y���㳻�C(�L�<v`�����h[g�P��<�_K<�4��g�ƽ�H��*�<�B�u�t>���=A��!��R�<d��<3f
=��<��>yT>;���	���=^��=DN���v�=�3�=��1�j ���X�:G����+���>.������=��>�� ���=M�>{%����6���l��]b=V^~>,�=Hr������ �=J!�:9ӓ�d"�w�:>�Ě���=($>�;!���W��b>�-��s��ƹ*>��:Z���#>��<2�<�}�p��<Iy�;�7=u,�=�q���u���^����4>��=���%��Iƻz�=ُ=��r��M>.��>�JƼfwH����{��=e܍�>i���Ѫ=O�ݽ�%ݼ�,=�=<f��<X��=Da�<y��<��u�� $�D�4���h<$��=�yA=�&�<ٛʽ＞@��J�2>e�B=�kL>5_�<8������Y7���ὑّ�0��*��-q��Z2��̊ƽ\X�>��Ž�e�<�ɽ��w>\��=�oͽ�I�<w�=�y<��ݼa�8�F���b�P���=4��+:���%
���'>u}=��u�
��=TR6���>�ߎ�qK��ֽ�Џ>J�=KV�=@�>b<$�>m�=�м]1Y��� �0�(����W�>� ]�v�>s�`�'�=�e/�`j�.'����%��=�q�="��"O��Md<Gޠ=ɦ��&����FľHR>8��_o>��=4k'��LT=�л��u��fS��
";�p�<��(={;Bn��S�����S�����:-=�a�傌���&���>�=Rp=K�o>7/���� ��<5#��l�q>�>�=O��>/:����9>1¾��'���=��<����$>������!=x<���ѱ��M�x��<��Z�����Wnc=��<�>K褽9P�=V��<�o>xt�$�T�}xý�5�!�=t�R>��=� 5�<�^�=5� �.Η;���#�����.JĺSf�: +=,0>>M�)�==��9E�=�t�W��-ܽf��=>�P<��w���=�P#���8>Vs�=�U��":<J���l;Ǥ����<M�=]� >�5J>/){<�2�=G�����9��Ƚ�d>���~�����=��>��u>���;���<a"�=�g8���8=��/>���=g~�>Q��k�ܽR��!����< �߽B�=���=#gR�ǀ��w�E=�H[>g�G>�>&>vD>�L�=���C�>"��~Q�=@��=~�><-�UOf>`��=�:�-��j�M=�p�*L6>�0�=�"����Q��>{��=~jh=�&w��ԛ>������=�I���4>��>N�㽱jB>� >(�=��<�� �a�>�Ν9
2> ���;ݽy��=ؿ˽-]�=�Cx>�����-h+>�����3={��=�z�=P;A��=J�(�@]�͢���������T���a���=I �>��=m7ҽ0>i!A=���=ͱG�ƪ�<�Ϗ��O���i��^�:>��<p�=�ɽ�A�<�"�j��>�=�����Y��ԭ�=Jd�<��=Em�=��&���߽HOY��#��܎=+�'����<�H>@;��ܽW9�6����m�<e)�<�.��?X�C�R��M�=W��=�{�<����#�����'���2Di��`��ڽ\���i*>�'��˗<-�>6�>v�s��>p؍>��*>�F>�}�����=8&.>|X>�W���+�=SZ �C�G=�����=G��/3=�5=!TC�	H�%��=�F�	���_�=��n<L����2�+��BO=��*�M9�=�轐I���` ��3�ǒ���gP<?+^>�|�=��'>�LR����nmR���=\E$�*+}�IE������Kj>(���=���/�潧;���G�A=ģ�<�W���G���V
��t���H�s�����.n>b����_w���½/�r>}�R��C�=V6>��H<Qǭ�m���=5jx��j�<�V�<��NPO�}4��{�������$c>��n��'�<��ݼڣ�����=8T�SM=5�뽁Ǣ=a�>KU�j��=a1�{����_=1ͫ=e����`��GG�иi=��M>�I6=1�#���*�]��:vq,�E��=P�R�1��=6D����_��,v>xٽ)����uڽ�ab=�Z���;��BnT�r6�h�j=cxb=�l�;B4���o�g�ͽ7�<Y�=gS̽�y4��;�=y`�<�{�<�ҥ��J�=�;Ѽ8���<?�G>#ҟ��->���n>v-��ҕ���+=�\�;��r���F=�)q=�"p�^�t�)�Y=)����rl=���>��L��:N��@�=D�E=��|�ԁ�|��ң�����b�=Xv����<�V�&��=՗���y�=��^���@G�`�i=�ey�M�;�ˀ=ø6��G�=�(�<�;�=0�����<�	v��>B>�=��'>v	��|�R3<r>wu��T��=9�	>PI!����>�,�FP�=Џ�<�(��7��=`|>ޜ�=��㝲<�E齅�O>B��=�=�L�= g�=����m�=�D�O����$��?콍��=r�;>���=[~;=���=f���)�3>rl�=���=#��=	V��I6���K�:��9��Q�<�5=M�> .���=ك>�ڧ��Y���)T���<�#j�3��=s���l��'?��;��|�=[=%��ۙ=U�z��F>�Ԏ<j��;�4�����h�<f�I>U���g0�=�7�*�c�,��<�ŕ����=�3>}&�=��w�M�<>�(�ϻ=��iƽތ��X�=*�:�z >���=v�=uG �["8>�r>�Q�<�@=V�U����=�C]����>g�=Fe<�,�=�6�����;!Å=��=�L>ض����7�ي�<�넾ȁ>�罍�=������yһ�;=H!i=����k=D�{�J��=Qn�Q�����=Dі����=��S��TT��P�\U^�a%V<A������>�;�����>�nR���/>�>�=�����
�=�6��"��=<�Z�[�;��<q;ߵ�0�v�K���G�<>M�> <��%=+��=1������<qE�,M�w̞��NC=�8#���=��m=0>~=�^>��<^Ȥ�|<�����~\��=;� �=Q�>x�2>R�u=Jx8��p��f�=�8�yH�&��=���<�~��۩7�F��;#���U�F>�g;>Z�+>���<���=�Q=)$_�?T,=W��>�Kؽ���E�r>�gŽ�1=_*�����S��Ѥ�樢>�w���O)<���]��Sg�'e>��X��;\�<�X�+�M��N2���>�f������&4=j%E<xvV<�[�</c=x�ļ������=4�=�@J�a�G=���=_#�=l�B�e^">O�%>|��>/�=hX�����7�=H9�ȓ=oj,�=w*>A�<"�4>�㚽c�ӽ���=�#��N�*�?�ｕ��Sk���;>QP=ހ7������qg=�f'�r´=�}^�T�=Q�q���/=�h=%_�=v->��=�e�3�������>��<�)=>���=����(�=e��<��=փ��g?R>�p?>j8=�i�V�<�0>�a>�)=�=2�w�->} ��X��=K�>��%����=�e�=���� �=�f��i9�@�>���<!��=�V=��A= �>�&�
�=�=m����˹���̽��;��<�d֮<��߼�M��q�?;9�����>(��<G!������t�=}����.�v��<����@P��(��&�%��@��>����'�X>>��$>ʯ��;�=]�#=���=�}��y�'>k��W�$�W�<[0T=�x8��Fh��dl= e#>�����\���g��fb��A�����<�Z=��$�5>>�f�<G��<��zU/>��B��X^=/��eY;�5��  5�M��<����JN>a˞��.~=) ����=N l�PY�;��̽]㟽�=���>��d�3/�^�5>���%F��>�����]��ཽl���H>ɓ⽅�c���d>���<�ʽ;"�<�*��=p���.c�=Y�<�=j	=�����7�@����q�<�6�<0P��kܻ{#	��C��߼:T.=.@�� z�<T~/>|��=��=�t5= ��>I�>|4<Ƃ>ezd=.o<��t��L�<�$=�>��=�0�<0��>T�=�K�\m=3�/�@E��n���;�C�<���=�I��K��QY�<��=�(��i M�9N=vv�<��潉(��Ե��n�P���o�_~:=���=���sc�Y$�2��<Fܔ=�I]>1�l�h�6�0�0��@ż���H�ٽa9>{c��<?��>��I=��$>?>��潕B ��V��Eǋ=��=݆w���=r� =g��3�	��́<~bٽS�&���8>�r���}��=��D�Z�*>>kF>#Z6=��O��=�9�<ʆ���#�{�����ε�=g���j^=�93<_Y6�%n�p]�!�9���_>;M��`)��<���F̜=���������L��=����"��q+���,�4f=�N�9TF=�y�=�w���� >��">f@=�>��<gn�j�t< �C>Kؙ<d��>M�]��J�=����ǝ������Ԥ�Q5ڽ��0=q���U��@l��%P�=��+=�7�����RF�<!��=�:���a>�_ͽ�#<!6g�#��<3�=��>ԩ���9�>��G<%��=C�<�!~�p[��A�n<cE��q@��>��<�_>Ӄ����=�	!�g�滌�ʽ���?'Q�� >�m���%��8�<��=y����:�=�䅾$s���������=}G'��F �w>:����>T��<���jM���>�,������g�=M��y�:=v�:>A  �uh�=7�I��&(�x/S�or>ij-�B�>��>u��=@��>	�=m �J�����=Z�=
����`�<�5��Ϗ<��n�%�=V���|*�z!=CKy=��=e7�<�>����f��oCK>ˤԼwEf>|�:���p=���=�Ӝ=�����/<����o�;�|>0r9�t��=,7�=��=�&=o�w�^b"��=�Ϣ����=K}�={�'<Z��6\3>؇J���Q�޽	��<+S�=�=\��K\˽��=UO�=mݽMI>67]>]#
>�o��o���wi>���=�x,>kٽ������H`ܽ�F>,.v=�
��8>�2bx�Q"�:�>o��=�~Z=������
=T	|�=Y��g��o��7H����<>Y�=D~�=f2�;1�B>��WE��2�yA>�Q��Ϸ"��nϼ�B=���5�+���]-4��U���?J=簆>����m���W�1y�DR=+��=J���ӻ��M�E	���&>��=�@q��_����><��}�1�e�V�=r>�>�R>3��]�p�}l�b'.��=>�x�<db����0���=�N���S�<_������ǽy=���or�=@0.�:��=��4>��v���6>%��=
ս&Ô<Ӎ>]?p���=��;�K��Q�{��=�;]Zѽ1+~>��W><�=�?���<±���Y�8�j������Y�v�=I�z>���"��=�J�=��H	>�U��|ѽnK���r>5���w�b�ׅ�# ʼ<�3�Wډ��1�7׼�k���}=�K꼇��=ĥh=���=���=5b��Z">�>HT���V/�����=_Ѫ>a��&��;'8�mc�=plJ����=����!>Xw�<�"����<��N>!(�<�;��:Z��i�<��>>������=-N9�V+��lf><��=�8<��6�[� �G<>|��A���V��R=�8d=��D>A ;�v>�������=��>㌬=�=>ɢ�=�(��:fg�ڜH�*���:���LW��{��M�<�/�V���TM��m��Z��=���=�4=�(�<5����gἘ�<L)�>��>>��=ꍘ��<��=�2���%�T�к��=�jg>�I=58��F�+k�==9�=
c���$�>e !�$�>�Ѱ=��Q>qp�=�	/����=��&2��Ǒ>����"�9>��&��wv=�<o>"�ܺl�Y>U[�=@z�z��='a�(�y=�9
� ��<pa��9M��9>tu�=�̫����=��ݼ���>�M���)�>+��=��ռ�=�;k�<�
�=�DK���v>�G��WZ=�L��M]�?�>��=8;�����ܽ�&]=�X�=�2�O��<��>T�3�����$�%>���=d;����=�ܗ=��¼*�c>`ս�5"=1�C��C<ض��τ=�"'��!M�o��=��<����e	>?��sP�<XI�=�v	�XD�='\�=&8>�_�=�p�8B=7�=�+�=� ����:�n��]�=�|�����<��e� ��8Q�::���=eK���隽�7>Av=]��.�)�᭒��=�c=̶Z�n�������<TX>���=\CF��[��r�Xn�<�-���==#�`1�%b>ޚ�=%�þ���=T�=��=1(�?[� e��~=GԦ�����~\�1@-=W��Tϑ���8��zk=4�x�n>y%�<����h��%�=�ά��Ţ�t�=��ü� ����k�a�;j�=�ü�{*>��>O�=��>q]�=�U�=�μ?���I�}���Qk���+>��
�8�=��=���<�Y��ZG��iζ:���I<��4=
��=�ae=3=6�'�F=��J=�g1��[>0���y�<�H��J���胾Ƒ��	>�Bؼ�?z>��=���=��ս�('><�&=Ck�=EI�=��=�'=�B�h��u:a��?���a<�,��෽=C9�=��<Xkt�����=d��<D��=��]=�9�l�@>��U=�N�=��=�ӹ���g��\νd!�#;�g=��ͽ�a�����=1ĳ>��B<O���@\<҂�M0��V� >�~[>|�ƽڎ�<����8� >S8�=3�<>\Q=[�<�����Ԛ=�	c��$I���;�a^=ɨ4>����� �<�� ½8�>(+�<��>D�ۼ]탽��	�B�=lV�=���=H9��R����=;�͔��4�=�v�=�#����=O�S>I݈��>j*<s4L�_ü=���^ϼeG�=���h+��m�����"�@.����=ul�=�)�<l\"��>��=���<�zR= U���[潝}���⫽g]=�:>:�V=�$=B.>n�N>����n��o	��^=��<?���Qq</���T]s��H��@�>ͭ=�^0�������h�X'��"<��n����@�=�r|=�]A��2�iu9�E��=V����k�=_-$���[>	I�=7���?���i�<�ث=fD��S��wb���VX����*S�m|�=�P�c��
��9%���ٽ|f����f="�Y=��ʽ �W��f�C��=�\콏�,<�i"=�B��L�wv��"څ���>S�=Q3G>s����>�d>]�r<�R��k@����.��~��h1�0>�Ş_>��~Xٽ�ܽ�i;�|Z=�D=���<��J����* �=���<�VH>�P¾�9�=߳=e
J=�tN=%I�ͥ��=�5���Ȭ���`<��i=��=AH>��<�@�ќ��-��>�w4�.]*�<���1d:��=S4�=��=����1GM��䔽��[=o�~>p0������=�Yc���
>c|�<�&@�x�������=���<
���{=��>���=�%ν�u=��=�L=U �HR�=��:���n=9Z>�*>7�>>a�6=�ؾ=ϸӽ� �={����0�K����7��5�X=���g��G><�>���w�
>�\�>�@�=��G>��7����=��?�����@�q=(@>�O$���>[Z���h����<>|:���ۺL&4>[m��w�=MLҼ�Z��;>�EH=��=5���1G�� ����H<Kx=|�S<VE"��z���wK>�(�=�׌=5�5����2��;h)�q}q(hhh(KK@KKtq hh	h
hh�ub�+3�460n˷~/��8�i�y�����;zZ�    iHJ��g���:6    ���/uy6I�6�:6T,�5��k5    ���UV��36%B6P�7�(6�f
�    ��K�nZ��y63����n��W�5zH�7J�)5�r�6�X糜�6p�7^�76:�d��#�>T�3�>�LK��Ӓ��>�2&K5�&�5�����6o�ܑ���4׹�    ��϶    ��5��6-�6    h)�q!}q"(hhhK@K@�q#hh	h
hh�ubEԼ�p��!et���R������>!C����<ՓK>|V����|�>�<�F�>m!>.�=���=�Y=T����$��E2<z0,=�S>��6�>��>O�q���
>]K�=v����=���=���Z�<b꾽���n��l��<>L�	�Fk���3=��>,�>��=��:>{@>V	���w�=��:Io	����ZU��i�>�ޜ=��t�&S�>����Y�@���FE��׾����о��m��st�=ٌr��07��C�>6TI���)>\���8�=cJ�<��=2�c>mM ;du��i�=l�c��R<�s$�����~�����<�p��c,�q�2>��Gh��0��� �p�5_���˽��2���д�<�ґ�G�*���^=�r�=�l����<P�>e>M�Y5�=�c龥H����>BTܼaz=ܯ=�L�U>$|o�P���=#��=*=��>RaH=Q�>�r�<�!>��>u4m=�6�=8D�<%���FU�=�c���߻=�f	�!?�=�~"��Y>����,�=����p�B=�>����<�y�=�=2�Q���=��,>�2�>�F>,��<�ߝ>{a��7�	>�|=��̾.�=>Zy>�Q�=q�#�\>�˜>��Y��b�h�K�
�X>z�`��$,���>+΅�jH"<�h>�s����>JU>F�8�ڢ���=|&�W�>>p��>!�\��RU>Oc$<سR>�3�����ۏ�!U*>&D>_!ٽҶ��9�>�\)>��57{=�Q}>�#�>�|��ۡ+�y	:����@/�=��F�e\r<����uM�>�r!>�ҋ>��<-��"��=L\:>�E𾌿�=���q�L������3>qD�<`vm=%��>�+6�*�h��y=-��=v2���[��6��]�+>�x�V�<=
zu<�*�=:�����ő���8>&�P���>�b=M�=�9(>��	���
>��h��=
��&b�=f��!Ľ#%;ӣ(>����V/�E�����<�ʻ<@e������M"�9���I�>I٤����c�7��ۼճ�>��C=�����=��<�L�=����@����.�a3>A�Y�i=p?y>��%�>l���FVT>������ܽ䣨;Vᚾ�s�=�,�=땟�Z��>"�R�����R���"�Ƚ���<��>�f�r�彫Z<���aC��*�]>=bE���=z%>Pb��ό>)��ý���$!�,��e0���ȯ=d�㾸�H�8���{�ȯ�=Z_"��}L>!ع>�WP���ؽW"�<{x[�/7�=��ֽH��>hҌ�9V��V���uv>�Ͼ���=��;��i=1�o=���������=?8�>�����<���U>��K��"�4O_�A�9�j�<>c��yR3>|\��vl�z.>\)�
�=�:��?��=d�=�RX=�*�= �=�
s>cg̽�-�>/.�=OLw>wX?��Մ=f�սČ��ѽ��=L��=q���Wh�����+�>D�/>`��=aU��W3>�4`>�V򻩮�>d�=S����仚�m	�>Bx-�� >�q�*�)>����Q5=~�>K2�oE�=nFS�7��<aG>���=�SƾY9>��{��@>�������|Y=1ɉ>�#�2s�==p^=M���CJ{>)Y���W����z-����>;r�]s�>9�=��ý<��<��C>B񗾇�g��ɽdk����������#���a�p�F�_�>�g=d3����>(���Ƚ6��J��J��N��t�8>J�:>��G>f�p�u�r�&.t>/G<�}:� E�;��,><~=OZ#>�A��P�_��x�<���=&E��a฾#��<�.X>��d�屯>5����>��%�����\��!`��{�p�>K��=�����=�Z~=+�V>�#�;���=Cܒ���#�-o�:b��=�~��։���Q�1ͺ�N��ҁV�֞ӽT��>cL�L��f!�p᥽�l<��e�.+վ�6N>q�R���P��]>���= +?>�@��{�ؽ_+���Fo=�Gq<��=���a�a�}�=BV�>�M ��1g��C�>�����ް=/�\>�j,���A��D�<1�=\L��ʟ(��z���<����`��
m=Lg����_������K�>v��=V��>�w��_�;�X:sL½!����ӽD�v���E>Yf>�X*���,>�4�=\w���Dp�+(3���<L��=��b>�%Z��NJ=�)�>��>#����e��P�n>%3=���<������<��F���6�Y|�;�>N�*>;��=�
����6���.>3)�A�>�y���T�>S��=��]���+���<h���{��o�>��'����= :}>��m='���o���޽��c>�ʽ�"8>6W@��D���;y��f��<Y<Gk��L{e��3�a��<�-��=j�`��>�F=B����@=O��<�ͦ���>�yz> ,u;1�!>������=�Ǽ:����>XX�=��x��?����j=#���`��z!>ES=V��<E�>4�)=��3� ��ּ>�{�>4��=�� >�>�=򙡾Ċ �
��ڍ`>��H>�٬� �	��`��<w\�>U�; �>���#>v�>��=~O>D1���o>�~=�;Ȼ��U=��	>��J>	�=���>ﬓ�K�v=*.��1h����&�u���Sa�Ȟ�=S
�<#�=0��=}>+ؽH������=C�H��>��E>����$�/2a��Ɍ>nd=zٽ'�=[Hj���ɼP�;(^i>�Q�>�~ҽͽq���e;s?u����=�_s��o�>&��>eʬ>	ز=}=����IbB=�f�دe=�,g>��>��K>z��=�+b���������b����<�	>P��<�Ǭ<���>甶>�:�>U��=T�j=�Y>xg8> �:ȅ���B^��'���ǽs�����>c��> �;���/7<M�O>�3�=�s2>��C��樽aC>-X>Q���"�˚�l�=,��s��-��$>�r�����>T�Ѽ��<�=�_ǽ�n���>A&*�Y��8�f>5_�=�� �J*�>�R�<��7>ƣJ�Z�����=���$z �c����Z��H�=}½iSa���=Hwj���d>Câ��˓��t����k=�J�>|�<)r�����d����>�C>.�,>�>�>o��Ծ<,�=Y�:>���>;\�)W��e�>��`�;�!�zXK>��<kۉ=^>��>��>�,=#H��	Z��e߷�q���`\*>c�(>��=��9�t��= >4��9F��E��=�w�=��>�>#���T�%�=]�'�� D>eꜽ�1�<0��>e5z�X>�=��B�m<-A�NZ�=u'��HϾ݊K�H(>T3>�Dͽ4K��0�"��+�=����a�E>{�v>�Y����>*������B�g=�g��o�;`�>�&t>dM =P��uc>)���Wd�>Ѵ�CX�=y�W�ڂ���y<wQ=a,=eG��ˌ�J��=h�9�\=��<�,��ޣ�=I��>.�{��g>ԓ�>=)=(����w{>u�������>�:t�o�;�ꤽ����>u䖾wL�=�SB>�����>֚��N�=�>�=�1:=�@=��ڽ�ؾ4�v=4�d�}s;<������>�p��Pֽ�����'>Z�Ƚ� z���̽��h��[��a��;���>~ȼ��+=Yk�p����M=en�=�����<���^���?=��,>i�>��7=��>c8<7��=��8&��U;�>s90>a��<*]1<[x�>ꌰ=����m��>�Q>6nA>���<RT�<훒�q��<J�ļ~Q"=�G+;K�?>�f���C=g�Z���C>�Q>�N� �=��=�ֽ"���FT�=[�'>��F�fڳ��G���׽k��<��2>`2�<���uF:��Fb�S��<Pݤ=qL=�� <�\�>���=k�D<���$ݕ�9\����?�c3>�Ҥ>O��>`�=>^>5�y>��$�[��>Pv='v;�T�i_c>����d�>���=;K���r����_�Q"�����9�=Ud��j>��<�E�=XXa�|?�[­��ؾ�^�A�|�HW¾�n�=��A>
d�ǁ>���=j�T>1�=$;>I��=��ψ3��A��t��g��r��>N��=��W�F�ܽ�z�<�u ��>���11R=)���]S=�v�=��پ�`�*���ݒ�GjC=��V�6&��k�=ב�=���;���=�R5>wtY��^=���1��w>�=�B>>���G$O<��}X�=M�½��>>Q�f>WPF=�\=�'�a��=�;����ǽ+O=*C������c%2=ܽ(S��5�-�\�׽��(>]7_��Q��y�3=��i�㐣� /���s>���>uaZ�<��=�'o>:^�=��J�`䬽��=���>u�=6TL>��*=�\F=8����M>��ӽ�Tv>�����h��?�ýu�5=��v=�hʾZ�A��b����n��[��-�=K�y>:�>�R�>�3>:pg>)���y�=�+t=Rð;�$��u-Q>�����fD��r��X��<_yq�~��=z���O�O�eN��5�a�2�47]>)/�k�>�����=�\�>-����(=������=�q����=�J>]�����(�J�y��:d�s>���=g=���=�f���X�>hK��_	�<�9���>�� �cz>����C0ξ�ڴ>W��=G��N@=+��=l�_=
oX>	�=a���y�=3Ë>!��꫕���,>�V�>
߼�B��z�<�&�8ǎ>�l��iss�a�B�Ӛ��tk�OH���A1��\\>��v�؈��e|�MKB<�b>l �����>ׁ>x�o��V����>��4>�@H�}��:�H�Qպ>,��=f��=W��;�V`=Iҧ�����C�>�c�<k��������>���'>8`Z�Q�_��h�� ��=9� >)��)�>���m��=	��)�=����l��:������=�|�;09�=j�6�~PŽtm">���=�=-Y�=��g�s���9�=H�<�m�Ļ�\��8z�>M�T�>�@�f���iX��n5>�V���F�=��>b�>���U�=���������c>�}�<�(�=Y������C�q=�nv>����C�S����=9��>,z�=���������=�ʾ$��_�սU�޽��̽�$q��~A>��J='�I>�U��
�=J����>x�0>5.>H�=k�a=�_ܽl����=uL�=�">i�=#
E�/n��c�=�����j;��=��=�ē>�tv��*���~�7�;�D��kŌ>�ވ>G�V;�����d<w޽�1>��=:�нq�S�1V�0�>��1HǽrԎ��}#>&v�>�	�g��=6�h>0��.\����<w�$���>�~�=������;�=t�O����~w�8�>1�=�>$>���L;3>%Ӻ�Do�>ŕ��l侘&���Y>���=���>���>�r&=ɭ�����9�>R!����=XDu>�:����=���K�\�W�>L}��ӥt<1�ռM��;X�ս�%D��*%>���0=�Ƒ��<�>,>��4�z���
?r`�������Y�C>Ah8����=���<�r���˾�M�Z��=lך=�MM=��8>�١��W>��/��C�����=L�� AF>}=�
�=��v�]�n%�=M)ټB�=�s��o*�`]���-�5�� ང�N<���\�E�<��=T�T>'�>>ћ>m�W=<Ӄ��0:;-�x>�>��>��=��2�=������5���a�V=��֐�=9h��='�O=�- =�V=xO��P�w=�?��T�=�tC>��>�����mS>��4=2��=�帽p�C�i�;������eb>�����m=�b�=*��>~ ҽ�Ľ�:�>J���>b���R<14�=A�>8�p>��:��Z<�v4>��S=W7]>ݳ��(���A���)>�'��g���:��f����{�_�n�y`��_fh�p3>8O����Oz�>͔$��ɽ�_����>p/-<UvO>ߚb�
�O�d��>25�<��������%���
=R��>�L<�#��J;)!>�*��-	>��<�!�p�ҽ�׹=��׽�yo��ܦ��˦>*?;��J>��^=F�x>�����W>a�>ϗ)>dZ�������"�q>�r���ž�9����=����=��3�/H>��l�)n
�1zؽZ?>f���R>��>�=f�d����=�`���f���
�>5/�>���Y<2�=�$�<���Ѓ�&�W=��>�,>]@W�6GF>2��>�Y��"������?>�F�>��>ݛ(>�2�X�۽!ɖ��r�>��ռ�Y�=���%>�=��*��
K:ݸ���=�^P�>{�=OS��R�>e�S���D>+����K>��=�Fp>�ya>���=�Q�<�[>�XO=�!�>��}<+�X�T�[>�U��T�>��=ꌲ��a>�X�M�=e
>m&>�Gѽ��J���`��p���y�=?7�>��*���վ0�F>i�춉��=A����>v�=�d��&5�'ؾ��ѽCP���+���3��m	="��<�������y��D>E�*=4ς>�4�b�T�6�?^d=��l>�<>u΄>S��=g�b�.���M�������Di�=�h�<t͌>ן��+�������B>\��=���є7>W��=�>5�X>3��铋=�"��7=v�b���5>��=��r�
N^>"~P�L���� �L ���Ώ>�hG�-�q��L�=��p��$P�!p�l�>��6�8��<tt�>v_Q�;f>�1=�򈾧�U��x���i��R"�^�=�Z�>����n(>�ؽ�����8=�,<h����*	�⋃���.��i�V6����=�V7;�����B>S�C�����}y�x�>j�K>�j��>D�!>K§�g�����������̤�����C�������=6|)=�K-�x�l���>��%�^�� I9>�*�(퓽��<�L>��� �D�E>TeW�(B�z:��F]�?;>�u�=��1��>�	�=����-9G����B�N>ັ��{�������=��>P�=M�k>�U�������F�BϾ���=� �>�t>xŉ�k�V>/����>/�<��O�>�l>�א<h_�=HK4>X<�������=[���s��ss&=򉽊�=%�=��>hx�>�`=-|I>��>|����>���=�^\��>����=�� �=:@����m==�
>Iym=!��O �sk=P,e�9����k�h�9��Z>��=8��=ȿ>�ֽً=	���[��>�_=<)����&=�ׂ=�II�����Xb����<帗=�D�P��𿥾�g�< �D:�z�<R�o>�m~>r�X��o���?��A��<VJ�GSF<˒<=4č=��a>��c�p�<>��?g��>uϋ��
>	����1>�e�=Ѕq<��n>n{ļ�>��^����=��>y`Z�7��D��=5�>���#Ň>^���Wgn<�m)�a�>���=̧]��O��l`��V��ة�U�>*���y��＾��+>1Ҙ���ľKS$=��_=b��<Q~>��j� �!�7��ȉ>Z�>!$`�o��<U���1f�=&��l���/C�v��;uܐ���=�1�>
���2���>l� ��(߽xS�1Kw>lt\�����=<E��=O��=-�%>���0�<'G�=",=>u��K��e��&�=��y����!�=��v�R�p=8���nQ����>1�[>����<�>}&>�C�#��=�=��Tܸ=N5M�|�>�fn�_�M��,��I>�%���=���򾽯�1=g�O��Xv��9�=��>�慽|�<<��=Y�*>mta�Z��J��;p���u�>S� �2�|>�s���p=w�=8=���V��@�>F�b>Rkc=DM�=��:��i+>/>�%�=ş�=�9F���s=�b� �T<{R�=��ľH<�L�9!��⇽�$4����=G�;>�훾6��.e�Ν��r>�q����9=���U%;���J��Y�=�S!=�FT���/=�H�=x��=u��ż=���>>�>�O�<�?>����V|�'�>7�}>O��;����"�>�7���%>s��=��p�p5�=��>���<P��bh7�� P>l;q�b;^>��_>G��q��=y`���;��I=���<�h_��E���>������7=�8��@�>9�=�І�X�E����>��=��>�����T>����<�D*��{+>nz�=&[�=��`>�f��'�>K%�=GG�	��=9sY�����>+��<B/ʼ&�	��Q�=7�t�D2k>~͎��RG>��m>z�d==�O>�>G�<+�f>��>���>y�L>)ꁾK>I���ޚ%�c����"�,&����<�����,�>r�<�s�Q��2�O�v��>�G��X�=c'��X�<�,<�#H>�`��C�9�c��P>���=�Ճ=~��A����5��uk�寽=��,����Q>׋��@���W���!�<�?a�R�>��6<�8$>#=�Z�Ճ>q�>
8�<k^ �Ls�=��y>cRR��=��A>�c>�^���p~>j��=�p�T��>��ǽ\~h��G@�������5<�[��e�ܽ�h���m�=aTf>
(>L*�=�����=�y齆�<m�M=��=��=d8��)��>~� >8��
Ŭ=�>�ō�O��,#�<��ս���,��Y>L��<E�=Px�>A��=1,Y>���e2�;j��16M>F���y^W>�2�>�4Q�R�X����_���:>����y;��F	�ԭ;>��Y>�:���>�E=�(�^!ȽX�=�G+>Ö罷�¾�<"=8T>�=��=�y�
>�����U������>���=IRo>�$Y>f�Y����(w>`��v9�=��∸�1�=�
�=2
 �j۾�p��:�>��������K>�����P�>oE]��d�%�O>�*#�����=+0½�z[���=�m�q�=���/=A�>����̿<'�ʼF\��2F�=M�I�G�}�*����O-Q>w���{��{�x=��e~B�%��=E�>�?d����=P�=��ۼ�r=��\>�kW=Ij>-�{>=Ph>���>���mVϽ�徻�>��>��Y�e�=�P�=8�@����� �m4�y��ۤ%=�3>;6u=���=�x<��<��=�u�=��D>�.=d5�=*}>R��=����0j9�3�t���>d�t>�)�>nS�>d�s�;=
O��j->�1��!�=�:��z��H>�]��6=�=�	u<�ϰ����Z�%�<=	�n�$��>&	����={��e �������f���s���d�=6�������-չ>�d��j׻���S_��yK�t  ��b��u�<!�>�ӽO��k_�8sʾm��k����J>��|�I�i<�l�>uG4>�D��	�X=��=�kx<}6��������A�=���/�=vp>�▾R�2���t>?H���6�=��%>��8����`��=���Y�����_>�*i�b�=�xz>�1��C郾x4��>�V�$�k��|���`�'=<"�>,ed���L>7��7���4�T�[�2<��ѼSW˽D�=c�>���=2?Ž~�>��A<�z�>eS��2D��p2�=�J�[�D>�W�<��l=��=�h��K��,�<>�>j��pZ,�5B�<A9�W��=�\S=�빽�vv�9�X>�/%=m=����9\-�\�>�o^>��:��X%�<x� <�b�=�.<�΍�J�w>�u>{>h�>�3�=�»�=�*[�ᇎ> ��N%'�MTj���=�>N���l*��*�H��>�"r���`=R�t>��
>�b�:]9����	��F���&�F��>�ȁ�2�?�M���#����=d�p>\�����<MH��r��{P�g�&��q�W�=8;�=���>�\>�	>Pء�8��5x���>O����`Ľ��	��+>
����*��MĽtժ=Ș>XB>���<� ξKhh="��=\iU���{Ľ�",>!�*;��I�1S��r��;0bm=�Ч�_��D�Խ��/	��z�<�9���0>��=�m�=sŞ�d�<PUb=��<�|���
=��_�R<�Ɨ+;Qb7>VO�=��=�w�=���ԛ4���>M�<>���=�,���=�K�����=y�<<�3�>?>{=B���Ȑ}��>�kT>@n�=a�L=�L>�C;^���T�>\�l>�WϽ��$=��I>��n��B>=4X>`}�>\.)>c�$��] �H&���J>ر�=� <�Z?R������=�t�;C�=�(�>��3�t�7>Z��|a�<Y��=��X��?���ep�
Jm=@��*p��=���>��>Vܮ�)�:>6��=H0�=}I/>��=�0q��m�>s�=��s>�k���+�<�I�=Yz�=����!&�z�����=�Q���$齁Z��$Nͽ�Rb���=s��>'H��~֍�D����@��U�����>�۾�M���^޽?����Z˼���=;=m2�=�M����[�����@>�r���;>3��%	��j>��<�Q���;�p��T���M>V�p�N=�o�=���`@>�i>W�;�.㌾��>�����>�l�=05�=^J/>�.�=��<�������~ƾ��!���=��k���ּ��={@�=�o�>��W�4�c��CZ����=��ӽH=�=lpH�,��>�<;(?�٠��r}��`{> �>��U=A�a���0>�g?�ߥ>���=��=e܇��?;�쪽��P>��8�<C��HT�	휾��>��<;��<�-�<ꨋ>�84>�>2�6��wZ><���=`8�=���=f�A>B͌��쀾&��>vC�=�,�xW�>���>U�k�+��=�EE���>�Y��Ip�]�]���>PW�=m�s=��<�ֽ�ZM�N�>�Q�H����q=�Z>��>,�Q��	>g�>9ڡ��!>�:�Av��FN�l�W=�۬�˯R>n��]�=���,��q��>����/؆�p7=��	�q=�8�&>�� >[�5���;>��c=��K���;<�Ⱦ��8>r��=n�R=3<�@�E^��=苼1�6>�5$>�:���#>�9>�S
�P;��^n��)">�#�5�P���'>�l�製k�;3���B���A뽽��r*�>�*�=�v]>��T=M�$�K�����>u�M;��¾mVt=���=��&��Z>�n]>2���iͷ	�>����Uds��6��ɝ�w���3yT=͜���;�:!<���ގ��a4����>�k>r�����Z=R� �F����=ٖ��O�=�����T�>	�=ʰ<�/V�{w>>8�s�Paq>(q>��ȼ�B��8w�<�2�<���=l��<OJ#>C�Q<|�A�%��;��� xi�-�N>� '�!�>��E�=`�Ț��.ꢽQ�>o���9���>��N>v��k� �>ߌ��=r>){�>��k�՗�,�D���>R.=r�2ػ��N�pY��)�=?\<=��>��>,��<�\�6��t&�ס½�{��Fq>;ļ� ���=��\�&Ve>�D뽚�������3�z�-���y��x>����A�z>H�J>�I�c|�>�ϔ=T馾c�R��������� ���=���==S�Ujs��Ÿ>����(!>��=��뽏r��G�����>���b5�>�����b�=�*���:�T��ǽ�C>CQ�=�=L>ǥ_�K�=�=[����X�����<�,�k4>�͙�#�'�d��;'N�5>�-����	G>(?�>�fA�b=�>H��<�ͻ�O��K A=�l>�O�����������l��=��<��_�Ȩ#>WF���<��>?�5>�b>x�?>r1>+S�<ci>oʽh�<d�׽?x���C���>��D=�\�=�>v��=��(��!@=�ӥ=��>ޠ�>db=S�����ǾLM>��3��X�=�'¾��=t����1�h�
���M��<��7*���XL=���>f��>��2>�Z8<O
�=�>�"D��A�<�����ۼ5��=l{�=�h�=&�?����=��V�n�3��=T��Q >��<��$>+~:���=+��<�^4�]�����x����~���Xc>}>�o�x��>�0��Fi=�h>��t>�V��@���'�t����p�='a����B��[��>�Ȋ���>V��e竾�u�<�t�<�b>��-=�Z��[=��<>nk>< >�0>�<�=�g���t��Y�<FR>P���W=ӽM=>.�[���۾uo�=y�'l�=q��VI��K������>6�;@��k6�1��<,н�u/<.����=���g>���=o�n��|>��>H�T�x����>).9>�`>�@��Z�=�f����N�=;�=|�=	~��_3>*�߼z	��A���{�=@�	>v��g\{�i��i>��ZrQ��k�����=�I6�&�<�>�[�<5IM>$�սb�þJU���=A:�=rI�+�=	d>�0��1I��t�܆d�z�P=�TR>u�C>�>���-0%�䍡��4p>O��>���=�n�>/!�<ǔϽ�8���2�'
����=���]>�-����=�#�;4�>>�T=��X}=�ݯ>����H���|�=5|l=|z��`����&����;7��=x�t�ta��9���>�>�һWb=��>~�K�@!.=��
�������.�=:Ծ�����P���ߺ���˄���5M�>������<
�?>!���	a0�������E>�E<��]����=�0>���=
�>6|��L�����U>�JŽ��^>��H�J	�=�>Ƭ}�?�?��ܳ�y�=�Z�>��=������j�ވ��F�>x[D>J�����=+�����3�%9/��l�=�r#�u��=!��=hx�>j�;|��v�W��0��ja�ɓQ>,Y�<!=�=hm?���!��X��k�p>vJ�=��>ojd>�~���~ �qD>��W�j���Ӽ��#���<'��OIh���>ꅽ���l�P�(=
B��	1g�~�%�v����yj�����o�c�mܫ�2��B�(>"�=�j�ٮ���-7��]����=��=">/�����?�Es9>c�=��Ž]�J>�.���c+�~B��S�>�>F;���8�h��=.�ѽ���g�=��Q>�~��HL>�6|>�����u�<OL�=U���O@� ����>W������>+ӆ�w�9�6&+�����O���37��H���ȼ<C>�sO�=��2���i>vG�4��=�KD�ǟ���GD�W�پލ><�Z=�T>��c���=��",;=~r5�R*r�ﲴ=i��=�I��j�W>P�=��E;��<�շ�e�����={B�X�"�\���5�S���� Ͻ�$�=����[���;R��b�=֋>Z-�>���H���D2����,=�L�;�̯>�]��YQ>�:@�%�!>e0�;(����S� ��,>��=2�=�ۓ<@���N�t>|ty=Y��=�Y�>oy>���=[�S��Ґ=6U>/��=���(e ��ָ�M��������=j�>Q0�>:Ɯ�B�v<�x���]>J��>4>C�����>:�x�����¶�f���v�<�%���}����<�J">�$-�[�=�w8�]�J>$bP>���=��/�F��=[��<���3G>gH�<֗�R���#����0@��v!�YV��V���[�v���X��>i��=d�:��
b=ŅX�g�;�	����8>Vs=�<�P�䨼�T��+����O�`ž��-���Q>�ƽ�d��v.�i�=�z<�Y'>]�=ZP��P�>�}���X>�=lͻGج<��>я>9���Z>�M|���1;�yx=�EZ�i��>JuX=WOI>1��Ǿ���=��C=2�h����>�L���2��b��I���c���w=�J�<�Ƽqf�<Kw=J�<���==��=�H>kg�i��=�J�<�5f�5��>ZĬ=�>
Do>~�>Z`,=�p�=�L+�"���������W���	��V�>��6���.�*���+���)��sv��@X,�D�>qwe>`*;>� >τE�[
^>ȳ����g>���<a���v�=!��=��w=�v���鳽N�$��g�SU�>�3����=������:�>��B>��ʻ�h/>=o���
>�P�>R��ˍ�=_�y<��">L~�=�u7��3/��k*�l�ƾ��]���֨>n��=��<V�Ľ'L�}ְ���d>P;���J�=U��<�ۄ=�K�>U{!�/-
>ڃ���;pr� �ھ� ���@��ܽ_�;���ua�1�=�{>�0��$�.7����u�I6)=(�b =K�V>ƫ˽n0=z��=��>/�=�!�c�˪�v�<CR����>�=7�\>��r�����V/>���<�����!��B_�;�E�>�ܽM��:��t�	>C#M��ַ��<�=>L��2ԼY7��Ȫt����>�l>f1��F{�=C�=�r^��e�=�p��Б�{�=�=$���3\> Y��{�>� �����=S:�F��;�m�> $�v����=3�>%2�����M��>V���B$p>�Ҕ��<�?>���=��>�����>E�x`��&�$��t=�����=��@���>t�yϪ�A�c�A~�9��>v.��/G�*�w=�6~��['�sƽڒ4���;��.��W�=G�7>��n>S�0����>*vý�������/->�J�>��<p�X=�_�>��4>C�4>�|1�/t>&.>B�x>��<6�;�a���K���?���;��=�6l>Y��=8'�=(�3>)��<�� >�q�0�ǭ>[h����C��ʼ��ս[��<Y�>�6>�S*=uȦ��/}��,��9ƒ�Y��=��=z�>�jH�6B�]z�>q���7���An�vH{=k�;�@������E�����^Ր�P^`<���<��>�@>n���ꐽs���>A�K=r�>>T\";3n=u�=�>�Ӗ>�9>6o���7L��}�;�E���+��<�W�/>-~@;�!���3>�	n>P
��J���>�У=�X뽊��Y�o>�<,�:>ʼ��q��|��=B��=����dF3���>�BY>� ,>Zغ�g6�<�,>�R�=�@�p,�=��=F�F翽<��>�9��('I��=#�{�[��<�$K�,�[���^���?>�u���檽Ma�6��<���<�%���#a���(�j��=ԉ���}=��<Y��)�_�}ھ��\z>�9���>5֒;B5O���N�D����f>����â='&Q�?G��Y\>�n+������*�}�R�򦦽.>Z�3�� �k�p�+���-�O=�����d<=�q��Dڽ2�T�;ϸ���z>+����>��ӼL�=�:R>�\¾��0�#.2�҅<߬	>�o���/r��s{�FR�l��>kB��`�T������=�ꔾL	K�!��=��>g�9�,d�=-P��J=�a �ʕ=�k�Cw>�{�=d9�=�_��"^n>�<�H(>9m�>/�l�֋ｼD|�o�j�`��=*��.h>b��
9ʽZ�=�Ǐ�I�*�3>3JY>���=z��>�>��G�2>�߰�JX��_a4����>����/G�>&n��Ե���Y��h���Ҥ�v@��<R�>4��MG���<f�O���I=<;Rim>��=���>�h���!`C>`�t=��w�p�N>Z�v��+�lf�-�<x���^b-�ĿJ�����=%�2=��=����F�^>���<a�q>��h>�᫾�PJ���d>{�0��1�u��>��=��>k>�G,��ސ>)�����۽�������U����=��׽�e���>=�V�=�n�=��V=� �=NE��@����'>�^��_���g>�`>:�+>Y͖>��3>W�>���Z�>�Q>�ѻ�j1侶�|>#UF>��S>r��=V��;ۥd>��>�i�=h)�q$}q%(hhhK@�q&hh	h
hh�ub@��22�K���E��{0�Q�����3h��عh3�'K���޲��31���ǈ�2)����w���b��?v��&�P��(�2�q#���e��\2ji3��3��}1B���XӉ����1C�9�F]�1�Iv����\^���93u��2bq�PR!�T7-���������F�2���d9 226>��7Բ�&��;2��`蝲�	������
F��?L3,*I2C��Ʒ�»T�L:Z3!��3��W$�7�93�k6�Lܞ�ޤ��h)�q'}q((hhhK@K@�q)hh	h
hh�ub���椾os��м��^���>ϣy����=�c�<HP$��==��׾��<xcֽ��Y�?_�M,9>L �=��i>#(����>���;�L�j��<@7�=~�=�9#�z�z;FM=�i>�=�>���)mټ�a�ü���x�=��<�"��8�>�W>��-����=i�=�ƾh
�"�׋�=bl�=�Ǣ=].g<�Xf��2���G�m�G��D�vܽD6�=�5��cE�;��K=��>�7��e�u���*�R��>X�=9�>�΍�-0>��>���f@�H�$�*��:p�<�~�=;�̽Inw=�����T�<�[Ӿ�b��b�1�\>\�-=h^ż��ɾ��f�Z��`Q=y4�>K1�Ւ�d~�=
�O>ٵ
=EB&�Rj:>�eۼS_+��f`������R=s�R�=c=�	�=�w�.
��ě��f>RĚ��-C��7 �^潾�7�R���&��C?�<�M��~�>zo>=�+{=�ը�)9�>�Lo��G=I 2>M����������|M>ݡ:�`i�������>�ۼ����#��[����4�y������Rؽ�2����ӽ��B�ϊ=�s�>[�>q������%p�=��n>�8t�Ⱥ�<�Ž��>i��=oݽ���=��S>2s>�����/�K�>�k�<�6�T׍�;�G>J��=6�>8ާ>������2?>K�A><�>F4ͽ��.>t��=;��=<U����s�}�Q>38�>��/���<^S�&K��]�=$���ʽi۽��B�=���==V�����>4�>�����N�;�u��q=4�� v>��:>�L'����z)U��'>+̐��(�=��<���f���Ʊ��6�W�=Q
�>G�����E��2�v�Ǎ-��$�aZl:2�K=k5��޾�����V^�'g��n�>�ڻ���=J�>����;������=2��<sD��v*���5>�G>�"+�7;5�O(���3��nN��d�;��ۼ��=Nv�	+B�`ž֝�>	�<�ֽ���=Y�=��=(a�;�<�=�z�=�"�>��=(-=�	ֽ�>>2C>��L];C��U���+��e½^�`��H�����ʲZ��\>Z?uN��=^�<���="$�<���Ϯ>l�c=d���� >��j�>�O�<Ȭ��>��@Mg>�M>s�W=�Jս���=4a>K^�=Z�3�������`>�yj��H>�D=���:���=2ɾ�I=�Y��Y��Bϙ��}��s�==㰅�/�x>E��<=��=h͵�9_�>�g/>ݘ�=�o.�ZI^>#�|�:�\��(z����q�>Ю�>ɚ��O��=(K>`�����x>��.<�j�=��C��j�k�g>)��>���>+Β�o=�u����>��L>x9�=��>L ��D:>> =����w�f��*���D��
#�<R��=8&����伌�d�:Hɽ��龚�)=q���=7���B>��r=?`7�p�D�}���g ����=2�ڼ�o<�ｹ�>{��>���,M�����>�]�W��<l>��ｨ��<���=*VӽGI�>vׯ=��=Ů�=�ma=�?[��A�=c������!�oѧ�/�>l����8��0�z��iI<%Fj�4F>�e�>��&�Wvc��(&>̏�>N�'�=��]=�濽 ��=���Dg��/>N�8��+�=��n e=�Ľ�G�A��<?���b�<�9̬�ڝ�/�-��u'��*ڽ���=<��>N۽��</�;��޽N��=�=��qJ=^7>�|�W(>r�I>e�F��^�<�>�,X>�^>�"����9��a/��?���<�=�"ݽ"}�>�M�>�� ��!���5�<�Ԉ��F>�,��°B>*됾0�=���`=�=>���=,�=p�Y��8��JeںV�=Pb�\,�>����8�=$���	�>lR�>S��:�$��D�ѾS^�=�ʛ=Ї�=�]B�r��k����=e���tƽ[$�3�f��6>e�O>p�*D���N>�*!>j��9���)c�<Py�>@C���F>��>f�>�w�w�D>���>q�p>���<�|"�P�M>����=.Z�.��V�>��>%?�=\F���l*��l> �a�G�G>1u�>
j��E���7��촽�2�=�Z:>5%]�Z8G>(@�@��=&�= d�>�^��>L
d�@=���dy'<�>�=L1>F��='-��j=��5���=�j�=ۆD>�H\>�<���a��ɹA�<�M>H��۽<#W����;�P�>+}���=���=�O=�	�<̬>���A>@9=�����;_�@b��-���ؾ����l�$>r~����1>`�ɽ;�>pV>��?�`L�1q�>�"���s�>�~ؽ"%ֽ�4���+-�	j=� !���-}A=�;R=�m�=G<쎟<��H>�#9>�=��Ǐ� X��u^�>�s�Iy�:�y>� >X��=�[�p=q�{>{Ӽ�>U�¾l�`>��=�=����I>��Q=���>�$=eiF>�*.�'3=� ���^>q:�Nn%�X�#>��=R/���;�=�>>��=_F�9H���V=��=�==��������=8!��q��}>�{���k��r>�kG<����`޽��h>>o�>��7��
�����T�=]�=h�>e<w��3k��;+�-ۏ��%f��C��ٽ���=`"��%"c=���>�$�<�&|�*l�=�P
>sjv�{�j�(Ɇ>���=ƜƼ�䀽��5��J�9~��Bl���뗾�v>��>2��,��%�~�U��=��:����=��š!�P�=���=��=yW�=�������=�,=2�p���������d����9>��޾��>
�
>ғ>̱�;��:}�;��4�Ē���>��X�������
��j\>dB�>�wI>B%�J��=P��|�>��T>�2_>�,�(y#>	y>�p%�y��;5�>��*���P���@>����y��ӼM1����=�v�<�uq>��<B��S�������� ��/���~n1�����-w��>m�½E�%>����/>I��=��#���;>a�%�
<.>*�;>Cc>69��M��><����G?>�����Hb����=��b>�;�=�#�>����T����<hχ�!ki>����Ȕ�<���=�y���w�@ǹ=6����Ǯ�W� =~tŽ�uV=��>S�0�;>�����/�6U�=o<��ѽ�7=�b�>]u=Ԍ��P2�+Y>^�'>�`=�R=�h$>���X�P>��=��>]u:�^Bj>i�-�9���AD8>�Y->�k�>��J���=�j'�<�)��#��O��=n>߄.=�m<�c'�(ʽ���ܭ�>��J<�B>���=g�>��<�ޭ�;wA�AѾ؋�4>=�,��|��_��iX�<�"<�Q�=17������Y0��K�:h�u�EؾR�w���9>|}��Ai4>�t��r�>��>����9?�jv����Q����;w�=��>�����3>UCi>܄�=0�6��6һ'�T���>T��>��'~=�L���+�>�ڋ��ȯ=2�>��{�oĽ�g�>$����=�>��0lo��J�=�A��.�=1�5=��>Б���<M�U>���C�$�9^��o�=�.4������&>	`����_> ;:XQ�����D�����=��ݼ�"����x?�<���<�9�kL�U���I�>�v<�5[P>�\�<��r�����=�>��޾i�=���=m��<����d�=���>���=��
<'�=*P��[�>c��>1�W>�.~>�f��6��=,3�>���=��欘=�q>`꽢��>��	��C��=X�d�n��;w�����뽟\>O���=�0>*BƼG�L>��{>Æ��D���=C��<�@ּcB�?�>W<��LO���=�py>��ݽ\5m>('2�L!ּ�*>�/����>�=�/$��=������w�
�x-=��>�
A��>z��z���`��I輪�ڽ�,E����>��o�[����=�͆=G:�=�� >l���EK>w�>.^�O�=�*�>>�L�<J�,�c���}>�ו<=DD>�_�0��<�?��s;�O>Wl���ً<9
�j�=zMQ�(�`��ݽ��"�Bg�>ڱa>�|�<IǾ�ׂ��N�;�(����;F-ּ��X>��1�Z�>�d>�¸� =��=��'<X􆽔�G>%zS>�+=�w�e�<� s�x�2>�\/=e*\���f�����CD'���9���>L���'�=$��=;_��8��>5�>D�X�4N*<�5��)�>Y�
>7��=H���۽o�򾱌�=�x��j�P9>W�ۻL���~F<ea)�����I1-��!.>B�l>�=�*�<�vB��$�=�K\��pM����>�mX���]<c+�NaA>�Ag>�@a���/�M���$2��9�=n"��<��=�u�=xw�՜��@㽭nJ=0��k��=��y���4��.|=S�6��g��Lc">p��:�>�W��2>DIͽ��������׌�GD�>��<O��>�=�R�����c�>��>̦���ߛ�b�<�z �z�0>� 8;$}ν����$|�x�軾�>�O>�j�=l04���E=���=1qE=��<��̽l�I�W��=�q�>a=X>�9�>��=>�Qͽ�86�C>>�d�u�H��>)y>�n�=om���@���ו��e>�P=�
>�T>JVm>~�����>��>��=�=^ᨽ�m:��=��X>r;<���>#C=����=�:=�=�鎼^o׻/e}>Ǒ>�a�=UQ����WA���p��o�(>Qv�=,b?=�1�>����/���8=��ҽ�\�=�z�=�0ҽ�ex�ҳ;=nO�>�%����\<���< `>=_>R��=��>��:������/��l�_��<�a>ո�=ۈ>����V<����н��^����=a��IQ�>�Nk>�ӽW�=��P=��罱��=<�>9��6����9=��3��\�>����k�=4�>*j�� �!r<cC>�Z��d�=Umֽ�~ļ�3�qʼ	k>�1�L9�<��w��=�[>��>��������!-��ui*>�>��<��u<��=%z���E������;�Ƞ����=7��>�z��۵� C��-<+;��v��:�>]4�����=�/:���8��t�Pi<�??>��|>����q+)��=b>)]��@e>���v��=�B��1�<*��>|��<��ٽ|-��5Q�@(ҽBq]=F����׽�iR��:�>EK�$�'>��=%m�����<�p>F��;�R�^ ���d=

>�=|>�	�lӪ��.���>0��0N�=��o��t�<	R�>�d�>V�.>ɬ��$�>|oZ����=�!==�6g=)C�=�!�=9�#>�
.;����&����A�z(f�kN;���U�>j=�@>c꽘]G�o��>k�B>-T>�ϴ>�Aۼ3���EY>�%���>��q�P!�/�[=�����&R����Rz>���П��r��=zL�<�L��Zt0�񟇾(�>��>ّ�<�n>Y�t����=]���%�>A��҂>�W���>6;�=����X�ߛ�;ˇ�=5_�0�;�K
e=4-U;��R>��*��?i=��M>�i������>��*>A��e-G��V�>�ƥ><��%��� =$��X=L�^> �>�є��Pn=ECQ��w>�<�>��1�|f��>!A>��= &m>�#o���B���g> �@�7 J>�4�D����(<r�T>?�¾����^�����=]b�=
a�>�WF�2�\>���=$�=ER�=FG{�Lى<� ��Qo�/[E>R�U�	|�=T����=!H���[=BTA>�U=�x&���.>V�=��̽G\�=�/�=q�3=Pz�>�����>>W�>�%s�����=:�>�~�������<"�s�n�9�O>��
��fv<
�ͼ1�=���=�#��j>��=�1x�&�=I!=P�#=�!�>���L9`�.:,>K�t�#H�;�O�����K���K��F�>F��Z�.��'�-!ԼW�=<�`��p>Gm�<_��=��<�����jM��`[>�v1�O��<H�>$��=ƈ�>���"d>E�:>a�$>�t�>�ľ�\���>�����1�_��=`�ݽ;L?Ց����=�1ս�U:�@=�WV<��<>�-�>� .>���:O �=��`���ŷ>�h»�l>�����=���=9@k>j޽nW=@D6<a҉���>I��=v�=i	i>����n ���ŉ�O��p9>�<	�����|">w{e�y�����z���_�%+�8�¾b�Κ�D��>���=�ig= ?����>E�B��4w�������9�_����.�;d���x�>�R�>���<��R=��ڽ/�=��=������p	[=g�^�`1��Nn>���=���=ߊ>l&t��9=��l��������<�W�A���~|�>����mS�=d��9�}>&>+}J>�=c��i'�={Bn�O�>I�"=��#�!�a>&�~�$�:q�#���л��=��<�m=QO<��ݎ�C\���>��/�"9=V�Z�O+V���C<=�=[�"�(���w�=�?7��K�:x>|ߑ<����v�&�ۼ�>��:��>A<a=�+J>����� >Dq>h�V>����A�/��:�>��!��h������q��)��@�
��T>͡F�� ��kB�=;=�:�>Џ>Q�0>β�����*|�X��=����o�<��=��,�	��=V1=�d�{}">1R�>VK���K�}�=Z�*���V>UPE�#2���~���=|�,>�Q�s��>�|�=҇�>�T4�|�×�5��<�-��0a�LO��[qT��?��ӗ�������<����T��`��>��:����=ij*�ܣ>�j
=�K=C�>���<�ͼ�e:��Š>2�2>����I=u=i4�>�����������!�=����l�G>��=f�{=��ؽɕ�>z�v��Jg=���EO�=��=W������-�=3~�7��=�>�o�����',^>��O�&9�=?Q<�PN=JP���`�>m��f��t��>&R��֦>�8�kz�>��[=G� ���½�$!�9�����]W>;�<#f>Rh�c`<=/c��z >�"콢�7>Oݫ��Kz>H��	���Q>S��<�j���$>�e8�a�s���q>������W��I�>۰��ʜ�\{�̆��Lq����<Kq��� �$k&���>�q�=e����\>�*��f�� �=�u�H͊�Q7=&��>򴿽�
��U��>��=Y���,�=(J�=�E{>3�|���=,臽�N4��ب=����KZ>Uy�㎃=�$�=�Կ�h�ʾc5e>�\=\Wy>�Ɵ��N|>�S�<ā��~�=NH��8�>5������m�����;_����=���=6���Kx�>��4>5H9> 
��<�ɽ� �����Fe�=h��>����, �>7�>���i��t���R2%>�RȽq�����>=��=���>�M�>�5ӽjǑ=�y�=
��g�>�O#>��>��b�`���([>��[�I�G>�`�;��<�bv=�����	�M5�=�s��5��N�����=�=�r7=��1�K>�?��<�<���;6c_�y�U;s�[>ǒ�rA���{��P��=�i�=����.Nn<6��<��=Ơa��L�>ͥ>?��_��=�ؑ��n[>�4�1��d;c��A�>���<J�=�U>��>�o<�?�=]�����4>�s��O���"�ۇ=B¼��<A��>��=g*:="ݽ�u">��q>^.��p!<m��M�= )�&Ba>��d=��~�I��=����U����R�>bL>扏������ʌ>�2>�#���M�=����C��Bg���=��w=ꉹ�d�=�%�9�==1�>]�=�+���'�w��=	Г�eN=�=5��������>x|�=p[�=�#�=_0^=����W�ݛɾ}s��*�;B�=�~>	k��q�H="Ʌ>�\�=�?�����:=��W=�wq>��=Ĺ�>k�>��>��=���=zs;>�b�=dRE>���b�(�!�>Ϭ*<��_�4>|�»=*?<��>:�:����1<>Q��>*>�<<ؼ�Ur*����>�YP>��<7��=1����Q�=oǳ�I����&E<��U=v�žT��!�ƾi���oľ���.��<�Sh>Ԝ��<� >��ؽS����d������c�>:Ɂ�).�r؋�t-2�0b�>��~�<9�ѽͿ
�"�Ƚ�6~=���Z�=+=��bư>An\���6�1&���Ͻx�w�h2=B�,��:���U����<��4��Y�=��>���9�=�{ �Ԡ�<^���۾RH=o�/*��$7�;�B�=�4��*K[;i�<��G<)=z�>X8
=�\=��ĬN��&��o]�=���6n�i4<���:�0��w�Sp�=�=>y��>qN�=e=k>��=0�0�׌,�_���=�C>�]e���>�w]>�L��C�n�P��>���=u)�<4Z���=>�/����ӽ	]�>�=�Md>�J>x�.���v>�� =Y���ç��	%>�ȓ>��=R=��";�s�B>�I@>�r>Z�`��KĽ^b��>�޽�-Ƚs.�v�3>�N>�H>�Km���N��`�>|X��at��)w����=<c��ڱ><�Ž�f�u�>u�g�z����ԾD��=�&3���\'>>6�W�zU�����U�(PF>��<�;׾��ƾ�1<>U�<ڠ_�2b<����i=�=��T=@nL� /�=0q��S>�$�>E�¾IVm�PIl=,r�=�Y-��pA> ��Q��H>9
��f� ���>_�ý/������=��=��Q�/�:4�>����H�;ED0>���K��=�i?�����}6>���3��<��	��E>�a>��4�d&��x�=j��=�b>�A#���D�6�<~ӽ��#>���>�ּp�ν��Gݲ=��=��^�X%9��I�>"��=!T�"���pd>[�Ͻ7�<aL>\_'��a^��qO�M�Q>rd��B>�
>g�T>������D$X=O�=�Г�����nI�PM>p]н�:��命��d����= �n>�����=�>�u-�u��=6->5����]���:��3m�H�/>P�T�'�G>�L= �+=G >�4=p�=3�w���h�׻�=���u|���>w�8���;T���e����>�ǉ�}/�����=N�	���,>��=M��=���=j�Z�(>@R��8��L4�4�>sQ=��;�� �>�=�O=9��=�gS>�ѕ>�ǿ=Ŋ�J���DнNe%��f���1ѽu���E�x��v#={'�=�� >)�=I�3�T��nHn=͖�L>a�s�[;�;80�~�=p�=
j��E�=���6O�� P�>�=�<�o�>���>��=O6?>ދ=�8�;���BW�>��>��k>�iF�]��=����@Ž��Òཤ�=�{�N;N>:1">9����@09vD���<zj=��(��2=f|｛�J>�(�N��s\���,��j-�=���n��Q
Rp��i�hh�<}J������c>��o<���-��~���O�=�.�譾���)� �h9��ȅ���=��;G>�=
�ԑ��R?�<��8=T�^=w�޽1*0=�e�>�B~�����=b<g%�=}up=]X�>�#Ƚ�W��0Y�<��>P��.R�k6��8��S�E�;I�<���;>D-���0���о��&>&9��ɵ|�����#	?�:��� �5>7�=���=�،=x-�������f��K�=���*������^����=&�>�ś��9��O=�fD>t>���>#*>��>���9|�>�kR�n�\�j	b>��4���p��^��/ݱ�bU�kB����R���N=>�\>�q;=��9p;f���Y=A�>V=4v;������k>�De������>=>b`��A�ɻ7l�=h6��*>)<�>��>�v@�'1˾לi���`��k�Eŀ�J�.�@�=�����͖�WR>�A�>\��y����<o'R�m���P(#��)�Y�Q=v
ؽ�%���R�<+��=
Le�@u��)d=��E�2>w�9�C�ڼ�W>�Ə;�ފ��| >5��k�=[_�gZ>���X��='s輻Y�=Za��H�>�������=�*��"���+�j�=��)7�����>KҽX�%��c�>��'��<Ōݽ:��i#ý6��yGq>�X��ٳ��S�%�>���}|>`�"��>N��=�eb�􀨼"q����=�l���y�����Ž���=�L���<[������m=�K¾��U���>�)��Ms���~|�ػ�Xr=�:=�|�=����D���논��̾�	��Y���2���B���N=�)�>�ľN��J,�z����{>"�����Jne=C~&����=����ֻ��=0�O�{�	>f�� n�>�=3!�>������x����=LM�;�Mr��c���pG����=�!>ݙ˼����8����"�jʽ�7k�'Y0��v��� >���=�ȼ.om�2�M><v��ƽ&�V>��½�l�=7�A�:�:��+=�۩��Cq>�L�=����>��=>Z�J������<`C:>A�2p>�:�>
?N>#k�����=��i>���g=����>фо�oy�ƿ���f���<��k�F)=��u>7U�>x�����C��k>}��>�j�=>�U=�q=�H%>%����Il���<(h��f��az�����=ey������>xM�=D~�>���=�
!=�p���ѽ��0�V�q>�B����=E3��	R;��]����)��/̼��<Α"�ٵ>~�`>��w���������K��Ԓ��n¾I�Խ������k������l�ν�Y���9=��;�Vg>"��<�8"�+{=1��>�Fr�?[�=��n=���=�e�� ��=��>i4>Elb="�P>��)>aU��[~���=ξ)R���n=2?��Ͳ��V�;yo�=K�Q�!���Z�==]���L�<��G>H�޾nC
=�!�>/Af=֌�=���=S��?�2>�ո�?��=��c�2|�=��=Z]�=;��L�����݅o>m��=k�l�\PY>l/M���>1��$=㹜<���H�9>�<����5�d�e�=b8i>w>���=R/དྷ*x=D�=�"���G�<L:<N�E���=.X�>K�>%�>� �>0�Ҿ�=>îǾx�<�i��r=㩽ӿB=�s���@r=~Fe�Ѭ�=�1=���=J<�<I'�=;az>^
<�u�2��Ž';��|h����F��7�>�=.K��z5>�+�*���1�D�k�П��6u�Ўؽ�`K>w{���X�>|�<�t�>K@G>&�|>Lx�=|M;d����"���8�hs> ¬=C�c=��%�Age>���g��KB(=O�=/��)��k��<8�=q�v�ub~>��׼K^\=�D>�����#=����Y�>��4>/=����A2*=����c�=]NA= [Y�"�ϼz8�=i�Ľ	�˽�Z��u��=ׅi=9�=V�*��ͼ1�6:�k[=s��>�Km>㙴�Ah>X~;s��^?����0>-XʽAѝ>�@��r��{�=�	a��nվ��m>.g��ϙ���3K>U[>�|t��]B=�N�=Kq�= ƾ>��>>l�ݽ�і>��>�U�>`�=�ϴ>! ��i��=._=�[>c2����Q��)�2��;�f=�I�=�޾4+>x�y��J�=�2����5�z�<�>>���+>����E���_>���o�$>>�@��a�R�=�Gʽ��=�cm>��R>���''>���=��<�9�NP�f����-q>N������� ����	�n� >��>}>y�Ͻ��7<1[���
��sv<4At�%/�>��=L���Q���}=��ڽ�R+>avI>�9����v>o?�>�6=� �����>�6�J���ʽ��A>�>»�5�>����C׼(�|>aut��L�>#O�=��Z�\�>tT׽|��;m>������:瘆�X�9��ٵ����=�=z��=-j>�|��{�^�=����Ё�!��<%� ��?����5�=n'>�������=e�>��<��,��f�7��>�^�>@��><����>RI���&
�ƊE�ƚl���޼wq����.=ڠ>=�=������>�@����}>*r�<ul��ٮ=Y�{>�>�IA>dm�@c�=Ǎ�=��N�g�=�{b��>}^=���=����x>91#=9a>�E��dÿ��cW>�|&>)\̽ٽڽX��=6�s�w���;?�<[;!=�`m>�tQ�$#�0z=$���|b>������>r���N1���B�%��7A!�c�K�a}f�_�ˋ�=c��=:E:�V����=J�/>S��8lX=Od6����=�m���J�=db�>�Q>N7�=:��"��=q�j=QDj��1{;�b~�.2�>�$���l׽>̎R�Wϙ��R����=ɨ2>���ԙZ�{ �=�Y���ql���O��<9*��4���jq�=H�>W:���}ʾ`�!�����TS�0���NF�t�=a�?��;ý莠=3R<_f0���:>����i>N
>������>�׼�"/>
�II�Qv�>F_��`�=�9>Z5p>g��i������#�l>�<�fv�=Ҁ.�i��˩�>�}�_)�:�Q��{=D��祺=F�!<�->��>�(=rT^�L?4�<2]�=�5W>�	�=��<��)��*Y�9����>,�W>��M>�h>P3=8��=t;�>�3��a >h�>Gcg=�ξg�C> b6���=���N��U��	!Z>�'��c�
�>��=��1>o���3佗�>>���>;3���=� �� ӽc5�=�P>�`�>����$5ǽ�#%��P)��=��B�J�｣v>��ϻj�!����=��<M>�w>��0����>��}�C���k�[���>��G�pL<����=<��>mʄ������=����5,>o{��|���w���ͼ�=�>^o׽��i��`��Rܼ�a�����u�>�M��?P�=��G>�{=��:��`v>P��=�y@���z�e&2��y��CL=�ʽPdE=�q�=&�>�t�� @���`=��c=1���Ž��������&�����=Ùy=a�j>s4"�f>������=[ּ���=�Q>�����0���;<��=VNѽ��=�dͽ�]>f)�q��Ɏ�=Wr��a��]�'�����@���0��=�6��I���>�i�=v��>�i�=�,g��>+�=^=���=?/�=_y/>
�Ӽ��D��^�=l�">�!X=�t>OV>;����X_>�/=�c3�Qel<f~w��W�<�`�=Q�`>�(཮0�������>����e}5;8��<�ٟ��p��cy>�>��u� p�>�g1>�����c>�?>
a��
����ν�Җ���S�c.�;�#=�U	�E\=W�b����������߾�k��6�*����=�[��nޡ<_����4����#<_�����-�/>��5�;白V�>�� >�쫽�,j�C��<aZ�>�ұ<8�9>���-���ϸ=��<.�\<3/u>�Q<��T'�މ�=�Qn<�H��w�<2�¾�¡>j$>V��0�>.�/<vU>:R> ��u��=D�~=�KL��2���#���H��ڼ|B�A��=`ڦ�A������ =X�#��o��;<~`�&��=x��������>��4���R�oc�=���F���e=[E����a=�l�=[��2��6�Z��!E>��ڽ�ý����ċ<�W��}��=K�Ͻ��=����q��,\�=3��>C2�>І�<<g=��>c�1>I�>w�:���q����=V�>>�3۽@�#�����@�2uU>�P>����K������<�$ʽ�+���l<�M�<kte>L�5>WB=��о�O�=�t��x/=��8�轒=�3P>�G�=�)�=g���cf���;�w�t>�q?�{���+�>0:ӽ��(>F.�?�N�폾�b��݈:Ԩ�>K�w=�">�&�X�>�pX>�<>"�#>l$��h�>yͻs����Z >����K=|�=�ч>2B���h>7�;�f������<�01/>���=	(���;0���j������>�^�����A
>��G�q.M�����>�s�>	<=1o½�བྷ�f�rB1���L>�$�-,>ȋ����=S=���-��F��>�½�a�}�<t�<����x�>�Y>����1,��(�=���DВ<��=�>zV,�4���p�>����/Y�G��>u�>�&��a��=�����o>U��=�l����K�S>'�p=�~L>KE使c=Y�����MB����3>~�>�˃>&�o<}x�=�I>������>�=�=��@W4>d[B�#�c�2�=��5ڽ#4������܄���^����=\�üq�%�N�����9�ފ�=��=�2%�b%��X��.N==�G>!�>�JG<�Q�=D��=ӂz>Ë"<齚;�\��O��i�*���?�c>�y���<���MSp>��<�;�=Q�F>T�%=�A��h�c>1�]��pc�F����6��y�>��V���>1����Х� .�=3�<Q���|n���<��&�N�)�t(�=�K�H+�=)���p��=x>�/%����=sB�;���<I>�>hͨ=L}��>;��%x4�`�%>э�����VI�{�M>�F�qj׼&�4�J�ӾP��@h>#��=@�=/{�'�m�x&��5@~;*��>_�}��	=o(�x�L=sz>�Rc=MOC>[��~^<lx����<�7��.`�T~�>^	>������a���;3��	0?>#R >�C���O���?>�� =��=�yI�Rq|���|�����n�����>@��=F�v=/;�=$D��B�=PT>��܁9���í����=:��=b� >�!g=��2�F�M>h���V>�#>"x ���&:#/K�k��%�=lj���4��p(=7c�bځ=b>�8��dI<�o�<��z��}��j�o=�B�=ŕ=��4>�=�>`��>ss��5T�Ьo�iҭ>g�\;sڕ���;�3���t��G�y��>��'�@�|=k5}�_�>B�V�؈Z>m��>z~T�&�->`򽊚�;,�3�/e>gA6�,F��l�=0g]=p�2>�1V=P��>]�I=�罅�½��>��= ��Q�=:�=y��;�f>�ꟼ`�㼲.-=�4Q��u��8�q�r�=�y5>B ��DN>A7+��{������Ƥ�>[jƽ�W���Bo>��>'��=�ٝ>߮���t�=��=��S>���=���>�~�=��.>�]��_gz=��*>�=��=�x�����>�{6>`=B���|>-� ����=�w̾,�>P��=i���p ����/��Ӹ��ЯM�)E� ��=�F>�.�����>B����=�{>��L���<l3���Ž�|���<m���5[��x�(�>��½�dq> ��I�<�^�f>{<�<aS����q��tX>�p�� ^>�K:>_{3=3Kj=�X�}����p�d!>��B�@��I�һ�!�>�yоv����1�zSh���>X�m�iҨ<P.�>ᡍ>���Aw���>�Rf=��ƽE��=%3�Y~>�r%������=��=qb�ġ���2>" �=z><��C^<g�3>M��0<����*A�L٩�͖4<*9F��¾L�,�>ƙ�/�=ҹW>�sm>o0��gE�����=�	p=��=����޶��6>�I>�Q��jo�>�2�=��P=��=mb�>lnFP�=�a< �׽�=#>N��>��<�d��$>�(ϽpJ�3���y=��<j	���� &��[Wq=�]����>�=��=5@B>�m[>������=�]@���۽/�ľDp+<{+!>�V?����e��>󨛻���n%t=���q�r��l=鯬�h)�q*}q+(hhhK@�q,hh	h
hh�ub�a�VT6����u�ju��܏5~��k�5v���y�P��6����U5N���0hb�.uR�������6}='6͸�5'�6m�6�X6UNM��{Q�'�����5��5��2�*��Dʯ4��&6I�ܵ���4�85�Q��:6џ�6v$S�:
�uA6�46��Y6L�˶$5uk��@�51�5��T6�0�6U��4�6<�o5
�Y�e���+[6TX�&i�����E���>6&6j/�6
��6h)�q-}q.(hhhK@K�q/hh	h
hh�uba-ν���=,�h�c�����R���v=?
�BLi=�qþ����`>ɢ�1�<#p��UB��v4��:���A�>�z>w�m=���=1�>��>�0�L�3��sŽ�"�=�K�=&��:Wr�x��<&>� ����<h�=�h3�0�>}>b5�����^�%>H>�:>8��R;=x·�_��=�˥=گ6>�>EZ�Mp>�}M=g;���н�;>�F9���u�ld����ھ�#>#l>
\�>�!`>h)�q0}q1(hhhK�q2hh	h
hh�ub�K�7h)�q3}q4(hhhK@K�q5hh	h
hh�ub�̚�9:��%�:���9�����:��m8�x!��o*:�B��}S�:j9��:��:n�:%���&�����3���Q��ʓ�?د���P�5.�:��:"���^!K�a���m�;����3 �E�n�yM�9ѿ92,V�w�X�#`�����:���9���:g@��)�8F�:��t:��I� �nO�8��:K�躝닺�K�栟:+ق�-U���M��y�:�n;����kr�W��98�:K�;ͼ������_;WL����>:����<49`�9%����;���:��k�Na: C�n4�i3:?��:�:�-_:���:b��:��%;Z�v9��:#��:����}�>�:e��:��:]�:���w��H9=��:XUº��@�9R�9�݁�Hh3�We�ݍø
n:�]4�����*�@�B�຋���:���8c��98�͹Ŧv��ZT��\�����_�B� |09����/��Q���s;� f�ɦ;������*�9�g;m������b���1�v9���ߛ��#9t����7�:��8��=�=�;��P��:���9�l��0�19f?]�Vv��7-]84�8���9[�:`�:��/�{���=:&�P9e�����,��V:��J��}�9�$�:t���;C:/ʹ�V�8-B�:n��8Vvʹ��H}���:��9�;6��9j9:v��:�o�����8w�T����c��8�	8�r���:W���b�ﺠ��7�l<9�������U)
:�'�:I߁�-�8�-:�J#�^J��� !;؈�:Ih�9
:�N��� ��w�ũ9��U
9w��:u�:���J-��ӕ:+]%:�[:e�T�:�:�>���;*�
���2�О:7�i���Aع%-���w�:	45�����K��:��2�۶��7:��:s��:Ϊ����jw�:�S�:��?:XW��1Һ�5��FEϹ�?J:�P��s?��a:NZ1�!��:�I����̺g�t:�nԺ�ɂ9�&�e�����(AU:���:��Y�;�����:��(:p䆹�:��l89V:���:"��8��u��B���~�$�-�8A|����:j9��o��:J�&��+�:��:�Ѻ� ݺy�_:��c:��@;��:��9�E�:���9U*�:N�8��:���:h�e:�];CQ��}x�~��9�`C���:����Wy�:)=:M���﹌K�ˈ�72���:��E9*'�:�:����4�8���9�/: ��88?�:W%;v}�7����\���ŭ9��f:�X��:;�س�����t�Dр�����7��|;�"-�r�<:�ݺ���������ź��'�6��>`$�M�?��Jc�\�
;i�T:l����úd��:m �����J
:V�:�OS����m�9���:�ә:f�^:a�M������C��"_�9k������:�.09+��8u�Q:�5�9��&�z�e:��9��:�p ;UK�:�*ɺ��� �:�6;CFӹ�[��@�99:�O:����k��);N��:�y;gO�
d:�@�8ȃº�n�r|�8̙�����ۋQ;�bI�I �9"G�FH��=�7�e'��D��=��lǌ:���:!�:�I8:u�:�\�:�";d%#�͞��\�:x6޺���:X�!;]"˺�y��50�T�90Q9�·�A,Ĺ�C��\�:��;�nv�9�,^:�:�93�K�O:�u�9��θ�����8��g46�
���f.B;�=":�̄�h)�q6}q7(hhhK�q8hh	h
hh�ub^���G�p�7�7��(�������e.